VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openram_demo
  CLASS BLOCK ;
  FOREIGN openram_demo ;
  ORIGIN 0.000 0.000 ;
  SIZE 1600.000 BY 1140.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 0.000 1314.130 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 360.440 1600.000 361.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1136.000 692.670 1140.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 659.640 1600.000 660.240 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1136.000 621.830 1140.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1081.240 1600.000 1081.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1136.000 737.750 1140.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 1136.000 576.750 1140.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 1136.000 647.590 1140.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 782.040 1600.000 782.640 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1136.000 286.950 1140.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 1136.000 1091.950 1140.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1136.000 605.730 1140.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1136.000 853.670 1140.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1136.000 13.250 1140.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 1136.000 1162.790 1140.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 1136.000 1027.550 1140.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 669.840 1600.000 670.440 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 1136.000 1523.430 1140.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 567.840 1600.000 568.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 1136.000 889.090 1140.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 241.440 1600.000 242.040 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 210.840 1600.000 211.440 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1136.000 1046.870 1140.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1136.000 711.990 1140.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1136.000 473.710 1140.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 248.240 1600.000 248.840 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1136.000 241.870 1140.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1136.000 267.630 1140.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1136.000 480.150 1140.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1136.000 1169.230 1140.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 316.240 1600.000 316.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1125.440 1600.000 1126.040 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 1136.000 393.210 1140.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1136.000 1062.970 1140.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 771.840 1600.000 772.440 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 948.640 1600.000 949.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1136.000 93.750 1140.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1136.000 409.310 1140.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 1136.000 296.610 1140.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1136.000 489.810 1140.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 1136.000 1275.490 1140.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 1136.000 1214.310 1140.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 1136.000 1549.190 1140.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 1136.000 373.890 1140.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1136.000 225.770 1140.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 1136.000 1513.770 1140.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1043.840 1600.000 1044.440 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 829.640 1600.000 830.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 61.240 1600.000 61.840 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 649.440 1600.000 650.040 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 996.240 1600.000 996.840 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 836.440 1600.000 837.040 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 1136.000 206.450 1140.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 1136.000 509.130 1140.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 520.240 1600.000 520.840 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 1136.000 1542.750 1140.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 975.840 1600.000 976.440 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 799.040 1600.000 799.640 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 1136.000 1584.610 1140.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 686.840 1600.000 687.440 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1136.000 499.470 1140.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 612.040 1600.000 612.640 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 1136.000 924.510 1140.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 1136.000 789.270 1140.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 1136.000 216.110 1140.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 306.040 1600.000 306.640 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 1136.000 1310.910 1140.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 455.640 1600.000 456.240 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 136.040 1600.000 136.640 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1136.000 834.350 1140.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1136.000 454.390 1140.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1023.440 1600.000 1024.040 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 622.240 1600.000 622.840 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 1136.000 976.030 1140.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 108.840 1600.000 109.440 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 1136.000 1204.650 1140.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 632.440 1600.000 633.040 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1136.000 1240.070 1140.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1136.000 782.830 1140.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 1136.000 1330.230 1140.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 584.840 1600.000 585.440 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1136.000 1153.130 1140.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 1136.000 303.050 1140.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 1136.000 357.790 1140.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 754.840 1600.000 755.440 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 333.240 1600.000 333.840 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 921.440 1600.000 922.040 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 1136.000 1269.050 1140.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1136.000 261.190 1140.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 482.840 1600.000 483.440 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 17.040 1600.000 17.640 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 867.040 1600.000 867.640 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 574.640 1600.000 575.240 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1136.000 728.090 1140.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1136.000 860.110 1140.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1136.000 29.350 1140.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 1136.000 1304.470 1140.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 1136.000 1558.850 1140.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 353.640 1600.000 354.240 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 380.840 1600.000 381.440 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 819.440 1600.000 820.040 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1136.000 683.010 1140.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 1136.000 1198.210 1140.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1136.000 251.530 1140.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 1136.000 1533.090 1140.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 6.840 1600.000 7.440 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 1136.000 1365.650 1140.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 1136.000 338.470 1140.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 81.640 1600.000 82.240 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1060.840 1600.000 1061.440 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1136.000 171.030 1140.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1136.000 798.930 1140.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 761.640 1600.000 762.240 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 295.840 1600.000 296.440 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 91.840 1600.000 92.440 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1136.000 570.310 1140.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 642.640 1600.000 643.240 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 856.840 1600.000 857.440 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 129.240 1600.000 129.840 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 173.440 1600.000 174.040 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 183.640 1600.000 184.240 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 1136.000 1375.310 1140.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1136.000 773.170 1140.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 734.440 1600.000 735.040 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1136.000 702.330 1140.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1136.000 550.990 1140.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1136.000 1021.110 1140.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 1136.000 277.290 1140.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 1136.000 84.090 1140.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 397.840 1600.000 398.440 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 1136.000 1497.670 1140.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1136.000 74.430 1140.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 258.440 1600.000 259.040 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 499.840 1600.000 500.440 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1136.000 544.550 1140.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1136.000 940.610 1140.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1136.000 1056.530 1140.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1136.000 1233.630 1140.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1136.000 1471.910 1140.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1136.000 808.590 1140.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 969.040 1600.000 969.640 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 54.440 1600.000 55.040 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 1136.000 464.050 1140.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 1136.000 1488.010 1140.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 986.040 1600.000 986.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 370.640 1600.000 371.240 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 435.240 1600.000 435.840 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1136.000 348.130 1140.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 0.000 1581.390 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1136.000 332.030 1140.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1098.240 1600.000 1098.840 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1136.000 1127.370 1140.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 268.640 1600.000 269.240 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 1136.000 992.130 1140.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 391.040 1600.000 391.640 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1136.000 154.930 1140.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1136.000 525.230 1140.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 1136.000 1011.450 1140.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 1136.000 1436.490 1140.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 1136.000 1320.570 1140.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 119.040 1600.000 119.640 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1136.000 753.850 1140.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 1136.000 657.250 1140.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1136.000 612.170 1140.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 0.000 1384.970 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 1136.000 1578.170 1140.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1136.000 718.430 1140.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 445.440 1600.000 446.040 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 408.040 1600.000 408.640 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 1136.000 1507.330 1140.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 1136.000 1285.150 1140.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 1136.000 895.530 1140.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1136.000 58.330 1140.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 493.040 1600.000 493.640 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 44.240 1600.000 44.840 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 1136.000 1462.250 1140.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1136.000 763.510 1140.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1136.000 180.690 1140.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1136.000 914.850 1140.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 34.040 1600.000 34.640 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1136.000 145.270 1140.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1136.000 534.890 1140.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 1136.000 438.290 1140.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 465.840 1600.000 466.440 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1136.000 985.690 1140.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 1136.000 950.270 1140.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1136.000 959.930 1140.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 1136.000 1391.410 1140.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1136.000 676.570 1140.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1136.000 818.250 1140.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1136.000 367.450 1140.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 1136.000 1355.990 1140.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1118.640 1600.000 1119.240 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1136.000 39.010 1140.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 1136.000 1381.750 1140.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 547.440 1600.000 548.040 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1136.000 869.770 1140.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 1136.000 1568.510 1140.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 530.440 1600.000 531.040 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 1136.000 1133.810 1140.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 1136.000 1294.810 1140.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 809.240 1600.000 809.840 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 1136.000 1037.210 1140.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1071.040 1600.000 1071.640 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 285.640 1600.000 286.240 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 537.240 1600.000 537.840 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 904.440 1600.000 905.040 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 98.640 1600.000 99.240 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 707.240 1600.000 707.840 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 0.000 1591.050 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1050.640 1600.000 1051.240 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 323.040 1600.000 323.640 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 1136.000 1426.830 1140.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 510.040 1600.000 510.640 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 1136.000 1594.270 1140.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 1136.000 1442.930 1140.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1136.000 631.490 1140.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 1136.000 402.870 1140.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 193.840 1600.000 194.440 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 557.640 1600.000 558.240 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 884.040 1600.000 884.640 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 1136.000 1478.350 1140.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1136.000 64.770 1140.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 1136.000 312.710 1140.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1136.000 48.670 1140.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 166.640 1600.000 167.240 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 894.240 1600.000 894.840 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1136.000 879.430 1140.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1136.000 666.910 1140.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1033.640 1600.000 1034.240 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 1136.000 586.410 1140.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 873.840 1600.000 874.440 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 1136.000 1188.550 1140.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1136.000 161.370 1140.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 1136.000 1339.890 1140.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 1136.000 1407.510 1140.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 1136.000 1417.170 1140.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1136.000 966.370 1140.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 27.240 1600.000 27.840 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1136.000 196.790 1140.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 1136.000 930.950 1140.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1136.000 3.590 1140.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 717.440 1600.000 718.040 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1013.240 1600.000 1013.840 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 938.440 1600.000 939.040 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1136.000 747.410 1140.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 744.640 1600.000 745.240 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 71.440 1600.000 72.040 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 1136.000 641.150 1140.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1136.000 129.170 1140.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 931.640 1600.000 932.240 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 1136.000 232.210 1140.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 1136.000 1082.290 1140.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1136.000 190.350 1140.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1136.000 322.370 1140.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 507.260 222.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 507.260 322.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 507.260 422.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 507.260 522.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 507.260 622.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 507.260 922.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 507.260 1022.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 507.260 1122.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 507.260 1222.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 507.260 1322.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 1027.260 222.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 1027.260 322.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 1027.260 422.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 1027.260 522.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 1027.260 622.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 1027.260 922.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 1027.260 1022.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 1027.260 1122.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 1027.260 1222.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 1027.260 1322.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.040 10.640 1422.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1521.040 10.640 1522.640 1129.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 90.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 507.260 272.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 507.260 372.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 507.260 472.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 507.260 572.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 507.260 672.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 507.260 972.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 507.260 1072.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 507.260 1172.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 507.260 1272.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 507.260 1372.640 610.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 1027.260 272.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 1027.260 372.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 1027.260 472.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 1027.260 572.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 1027.260 672.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 1027.260 972.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 1027.260 1072.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 1027.260 1172.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 1027.260 1272.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 1027.260 1372.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.040 10.640 1472.640 1129.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.040 10.640 1572.640 1129.040 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 156.440 1600.000 157.040 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1136.000 109.850 1140.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1136.000 824.690 1140.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1136.000 515.570 1140.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1006.440 1600.000 1007.040 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 911.240 1600.000 911.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 343.440 1600.000 344.040 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 1136.000 844.010 1140.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 1136.000 1259.390 1140.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 204.040 1600.000 204.640 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1136.000 100.190 1140.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1136.000 428.630 1140.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 724.240 1600.000 724.840 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 1136.000 1452.590 1140.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1136.000 1098.390 1140.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 472.640 1600.000 473.240 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1136.000 1072.630 1140.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 231.240 1600.000 231.840 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 1136.000 444.730 1140.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1135.640 1600.000 1136.240 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 595.040 1600.000 595.640 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1136.000 1001.790 1140.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 1136.000 1346.330 1140.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1136.000 119.510 1140.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 697.040 1600.000 697.640 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 1136.000 1401.070 1140.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 958.840 1600.000 959.440 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 278.840 1600.000 279.440 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1136.000 1249.730 1140.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1136.000 418.970 1140.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 680.040 1600.000 680.640 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 221.040 1600.000 221.640 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 418.240 1600.000 418.840 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 1136.000 1223.970 1140.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1088.040 1600.000 1088.640 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 605.240 1600.000 605.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 1108.440 1600.000 1109.040 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1136.000 1178.890 1140.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 0.000 1536.310 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1136.000 560.650 1140.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 1136.000 905.190 1140.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 1136.000 596.070 1140.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 1136.000 1143.470 1140.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 146.240 1600.000 146.840 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 846.640 1600.000 847.240 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 792.240 1600.000 792.840 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 1136.000 1117.710 1140.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1136.000 1108.050 1140.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1136.000 135.610 1140.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1136.000 383.550 1140.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1136.000 22.910 1140.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 428.440 1600.000 429.040 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1594.360 1128.885 ;
      LAYER met1 ;
        RECT 0.070 10.640 1594.360 1129.040 ;
      LAYER met2 ;
        RECT 0.100 1135.720 3.030 1136.690 ;
        RECT 3.870 1135.720 12.690 1136.690 ;
        RECT 13.530 1135.720 22.350 1136.690 ;
        RECT 23.190 1135.720 28.790 1136.690 ;
        RECT 29.630 1135.720 38.450 1136.690 ;
        RECT 39.290 1135.720 48.110 1136.690 ;
        RECT 48.950 1135.720 57.770 1136.690 ;
        RECT 58.610 1135.720 64.210 1136.690 ;
        RECT 65.050 1135.720 73.870 1136.690 ;
        RECT 74.710 1135.720 83.530 1136.690 ;
        RECT 84.370 1135.720 93.190 1136.690 ;
        RECT 94.030 1135.720 99.630 1136.690 ;
        RECT 100.470 1135.720 109.290 1136.690 ;
        RECT 110.130 1135.720 118.950 1136.690 ;
        RECT 119.790 1135.720 128.610 1136.690 ;
        RECT 129.450 1135.720 135.050 1136.690 ;
        RECT 135.890 1135.720 144.710 1136.690 ;
        RECT 145.550 1135.720 154.370 1136.690 ;
        RECT 155.210 1135.720 160.810 1136.690 ;
        RECT 161.650 1135.720 170.470 1136.690 ;
        RECT 171.310 1135.720 180.130 1136.690 ;
        RECT 180.970 1135.720 189.790 1136.690 ;
        RECT 190.630 1135.720 196.230 1136.690 ;
        RECT 197.070 1135.720 205.890 1136.690 ;
        RECT 206.730 1135.720 215.550 1136.690 ;
        RECT 216.390 1135.720 225.210 1136.690 ;
        RECT 226.050 1135.720 231.650 1136.690 ;
        RECT 232.490 1135.720 241.310 1136.690 ;
        RECT 242.150 1135.720 250.970 1136.690 ;
        RECT 251.810 1135.720 260.630 1136.690 ;
        RECT 261.470 1135.720 267.070 1136.690 ;
        RECT 267.910 1135.720 276.730 1136.690 ;
        RECT 277.570 1135.720 286.390 1136.690 ;
        RECT 287.230 1135.720 296.050 1136.690 ;
        RECT 296.890 1135.720 302.490 1136.690 ;
        RECT 303.330 1135.720 312.150 1136.690 ;
        RECT 312.990 1135.720 321.810 1136.690 ;
        RECT 322.650 1135.720 331.470 1136.690 ;
        RECT 332.310 1135.720 337.910 1136.690 ;
        RECT 338.750 1135.720 347.570 1136.690 ;
        RECT 348.410 1135.720 357.230 1136.690 ;
        RECT 358.070 1135.720 366.890 1136.690 ;
        RECT 367.730 1135.720 373.330 1136.690 ;
        RECT 374.170 1135.720 382.990 1136.690 ;
        RECT 383.830 1135.720 392.650 1136.690 ;
        RECT 393.490 1135.720 402.310 1136.690 ;
        RECT 403.150 1135.720 408.750 1136.690 ;
        RECT 409.590 1135.720 418.410 1136.690 ;
        RECT 419.250 1135.720 428.070 1136.690 ;
        RECT 428.910 1135.720 437.730 1136.690 ;
        RECT 438.570 1135.720 444.170 1136.690 ;
        RECT 445.010 1135.720 453.830 1136.690 ;
        RECT 454.670 1135.720 463.490 1136.690 ;
        RECT 464.330 1135.720 473.150 1136.690 ;
        RECT 473.990 1135.720 479.590 1136.690 ;
        RECT 480.430 1135.720 489.250 1136.690 ;
        RECT 490.090 1135.720 498.910 1136.690 ;
        RECT 499.750 1135.720 508.570 1136.690 ;
        RECT 509.410 1135.720 515.010 1136.690 ;
        RECT 515.850 1135.720 524.670 1136.690 ;
        RECT 525.510 1135.720 534.330 1136.690 ;
        RECT 535.170 1135.720 543.990 1136.690 ;
        RECT 544.830 1135.720 550.430 1136.690 ;
        RECT 551.270 1135.720 560.090 1136.690 ;
        RECT 560.930 1135.720 569.750 1136.690 ;
        RECT 570.590 1135.720 576.190 1136.690 ;
        RECT 577.030 1135.720 585.850 1136.690 ;
        RECT 586.690 1135.720 595.510 1136.690 ;
        RECT 596.350 1135.720 605.170 1136.690 ;
        RECT 606.010 1135.720 611.610 1136.690 ;
        RECT 612.450 1135.720 621.270 1136.690 ;
        RECT 622.110 1135.720 630.930 1136.690 ;
        RECT 631.770 1135.720 640.590 1136.690 ;
        RECT 641.430 1135.720 647.030 1136.690 ;
        RECT 647.870 1135.720 656.690 1136.690 ;
        RECT 657.530 1135.720 666.350 1136.690 ;
        RECT 667.190 1135.720 676.010 1136.690 ;
        RECT 676.850 1135.720 682.450 1136.690 ;
        RECT 683.290 1135.720 692.110 1136.690 ;
        RECT 692.950 1135.720 701.770 1136.690 ;
        RECT 702.610 1135.720 711.430 1136.690 ;
        RECT 712.270 1135.720 717.870 1136.690 ;
        RECT 718.710 1135.720 727.530 1136.690 ;
        RECT 728.370 1135.720 737.190 1136.690 ;
        RECT 738.030 1135.720 746.850 1136.690 ;
        RECT 747.690 1135.720 753.290 1136.690 ;
        RECT 754.130 1135.720 762.950 1136.690 ;
        RECT 763.790 1135.720 772.610 1136.690 ;
        RECT 773.450 1135.720 782.270 1136.690 ;
        RECT 783.110 1135.720 788.710 1136.690 ;
        RECT 789.550 1135.720 798.370 1136.690 ;
        RECT 799.210 1135.720 808.030 1136.690 ;
        RECT 808.870 1135.720 817.690 1136.690 ;
        RECT 818.530 1135.720 824.130 1136.690 ;
        RECT 824.970 1135.720 833.790 1136.690 ;
        RECT 834.630 1135.720 843.450 1136.690 ;
        RECT 844.290 1135.720 853.110 1136.690 ;
        RECT 853.950 1135.720 859.550 1136.690 ;
        RECT 860.390 1135.720 869.210 1136.690 ;
        RECT 870.050 1135.720 878.870 1136.690 ;
        RECT 879.710 1135.720 888.530 1136.690 ;
        RECT 889.370 1135.720 894.970 1136.690 ;
        RECT 895.810 1135.720 904.630 1136.690 ;
        RECT 905.470 1135.720 914.290 1136.690 ;
        RECT 915.130 1135.720 923.950 1136.690 ;
        RECT 924.790 1135.720 930.390 1136.690 ;
        RECT 931.230 1135.720 940.050 1136.690 ;
        RECT 940.890 1135.720 949.710 1136.690 ;
        RECT 950.550 1135.720 959.370 1136.690 ;
        RECT 960.210 1135.720 965.810 1136.690 ;
        RECT 966.650 1135.720 975.470 1136.690 ;
        RECT 976.310 1135.720 985.130 1136.690 ;
        RECT 985.970 1135.720 991.570 1136.690 ;
        RECT 992.410 1135.720 1001.230 1136.690 ;
        RECT 1002.070 1135.720 1010.890 1136.690 ;
        RECT 1011.730 1135.720 1020.550 1136.690 ;
        RECT 1021.390 1135.720 1026.990 1136.690 ;
        RECT 1027.830 1135.720 1036.650 1136.690 ;
        RECT 1037.490 1135.720 1046.310 1136.690 ;
        RECT 1047.150 1135.720 1055.970 1136.690 ;
        RECT 1056.810 1135.720 1062.410 1136.690 ;
        RECT 1063.250 1135.720 1072.070 1136.690 ;
        RECT 1072.910 1135.720 1081.730 1136.690 ;
        RECT 1082.570 1135.720 1091.390 1136.690 ;
        RECT 1092.230 1135.720 1097.830 1136.690 ;
        RECT 1098.670 1135.720 1107.490 1136.690 ;
        RECT 1108.330 1135.720 1117.150 1136.690 ;
        RECT 1117.990 1135.720 1126.810 1136.690 ;
        RECT 1127.650 1135.720 1133.250 1136.690 ;
        RECT 1134.090 1135.720 1142.910 1136.690 ;
        RECT 1143.750 1135.720 1152.570 1136.690 ;
        RECT 1153.410 1135.720 1162.230 1136.690 ;
        RECT 1163.070 1135.720 1168.670 1136.690 ;
        RECT 1169.510 1135.720 1178.330 1136.690 ;
        RECT 1179.170 1135.720 1187.990 1136.690 ;
        RECT 1188.830 1135.720 1197.650 1136.690 ;
        RECT 1198.490 1135.720 1204.090 1136.690 ;
        RECT 1204.930 1135.720 1213.750 1136.690 ;
        RECT 1214.590 1135.720 1223.410 1136.690 ;
        RECT 1224.250 1135.720 1233.070 1136.690 ;
        RECT 1233.910 1135.720 1239.510 1136.690 ;
        RECT 1240.350 1135.720 1249.170 1136.690 ;
        RECT 1250.010 1135.720 1258.830 1136.690 ;
        RECT 1259.670 1135.720 1268.490 1136.690 ;
        RECT 1269.330 1135.720 1274.930 1136.690 ;
        RECT 1275.770 1135.720 1284.590 1136.690 ;
        RECT 1285.430 1135.720 1294.250 1136.690 ;
        RECT 1295.090 1135.720 1303.910 1136.690 ;
        RECT 1304.750 1135.720 1310.350 1136.690 ;
        RECT 1311.190 1135.720 1320.010 1136.690 ;
        RECT 1320.850 1135.720 1329.670 1136.690 ;
        RECT 1330.510 1135.720 1339.330 1136.690 ;
        RECT 1340.170 1135.720 1345.770 1136.690 ;
        RECT 1346.610 1135.720 1355.430 1136.690 ;
        RECT 1356.270 1135.720 1365.090 1136.690 ;
        RECT 1365.930 1135.720 1374.750 1136.690 ;
        RECT 1375.590 1135.720 1381.190 1136.690 ;
        RECT 1382.030 1135.720 1390.850 1136.690 ;
        RECT 1391.690 1135.720 1400.510 1136.690 ;
        RECT 1401.350 1135.720 1406.950 1136.690 ;
        RECT 1407.790 1135.720 1416.610 1136.690 ;
        RECT 1417.450 1135.720 1426.270 1136.690 ;
        RECT 1427.110 1135.720 1435.930 1136.690 ;
        RECT 1436.770 1135.720 1442.370 1136.690 ;
        RECT 1443.210 1135.720 1452.030 1136.690 ;
        RECT 1452.870 1135.720 1461.690 1136.690 ;
        RECT 1462.530 1135.720 1471.350 1136.690 ;
        RECT 1472.190 1135.720 1477.790 1136.690 ;
        RECT 1478.630 1135.720 1487.450 1136.690 ;
        RECT 1488.290 1135.720 1497.110 1136.690 ;
        RECT 1497.950 1135.720 1506.770 1136.690 ;
        RECT 1507.610 1135.720 1513.210 1136.690 ;
        RECT 1514.050 1135.720 1522.870 1136.690 ;
        RECT 1523.710 1135.720 1532.530 1136.690 ;
        RECT 1533.370 1135.720 1542.190 1136.690 ;
        RECT 1543.030 1135.720 1548.630 1136.690 ;
        RECT 1549.470 1135.720 1558.290 1136.690 ;
        RECT 1559.130 1135.720 1567.950 1136.690 ;
        RECT 1568.790 1135.720 1577.610 1136.690 ;
        RECT 1578.450 1135.720 1584.050 1136.690 ;
        RECT 1584.890 1135.720 1590.130 1136.690 ;
        RECT 0.100 4.280 1590.130 1135.720 ;
        RECT 0.650 3.670 6.250 4.280 ;
        RECT 7.090 3.670 15.910 4.280 ;
        RECT 16.750 3.670 25.570 4.280 ;
        RECT 26.410 3.670 32.010 4.280 ;
        RECT 32.850 3.670 41.670 4.280 ;
        RECT 42.510 3.670 51.330 4.280 ;
        RECT 52.170 3.670 60.990 4.280 ;
        RECT 61.830 3.670 67.430 4.280 ;
        RECT 68.270 3.670 77.090 4.280 ;
        RECT 77.930 3.670 86.750 4.280 ;
        RECT 87.590 3.670 96.410 4.280 ;
        RECT 97.250 3.670 102.850 4.280 ;
        RECT 103.690 3.670 112.510 4.280 ;
        RECT 113.350 3.670 122.170 4.280 ;
        RECT 123.010 3.670 131.830 4.280 ;
        RECT 132.670 3.670 138.270 4.280 ;
        RECT 139.110 3.670 147.930 4.280 ;
        RECT 148.770 3.670 157.590 4.280 ;
        RECT 158.430 3.670 167.250 4.280 ;
        RECT 168.090 3.670 173.690 4.280 ;
        RECT 174.530 3.670 183.350 4.280 ;
        RECT 184.190 3.670 193.010 4.280 ;
        RECT 193.850 3.670 202.670 4.280 ;
        RECT 203.510 3.670 209.110 4.280 ;
        RECT 209.950 3.670 218.770 4.280 ;
        RECT 219.610 3.670 228.430 4.280 ;
        RECT 229.270 3.670 238.090 4.280 ;
        RECT 238.930 3.670 244.530 4.280 ;
        RECT 245.370 3.670 254.190 4.280 ;
        RECT 255.030 3.670 263.850 4.280 ;
        RECT 264.690 3.670 273.510 4.280 ;
        RECT 274.350 3.670 279.950 4.280 ;
        RECT 280.790 3.670 289.610 4.280 ;
        RECT 290.450 3.670 299.270 4.280 ;
        RECT 300.110 3.670 308.930 4.280 ;
        RECT 309.770 3.670 315.370 4.280 ;
        RECT 316.210 3.670 325.030 4.280 ;
        RECT 325.870 3.670 334.690 4.280 ;
        RECT 335.530 3.670 344.350 4.280 ;
        RECT 345.190 3.670 350.790 4.280 ;
        RECT 351.630 3.670 360.450 4.280 ;
        RECT 361.290 3.670 370.110 4.280 ;
        RECT 370.950 3.670 379.770 4.280 ;
        RECT 380.610 3.670 386.210 4.280 ;
        RECT 387.050 3.670 395.870 4.280 ;
        RECT 396.710 3.670 405.530 4.280 ;
        RECT 406.370 3.670 411.970 4.280 ;
        RECT 412.810 3.670 421.630 4.280 ;
        RECT 422.470 3.670 431.290 4.280 ;
        RECT 432.130 3.670 440.950 4.280 ;
        RECT 441.790 3.670 447.390 4.280 ;
        RECT 448.230 3.670 457.050 4.280 ;
        RECT 457.890 3.670 466.710 4.280 ;
        RECT 467.550 3.670 476.370 4.280 ;
        RECT 477.210 3.670 482.810 4.280 ;
        RECT 483.650 3.670 492.470 4.280 ;
        RECT 493.310 3.670 502.130 4.280 ;
        RECT 502.970 3.670 511.790 4.280 ;
        RECT 512.630 3.670 518.230 4.280 ;
        RECT 519.070 3.670 527.890 4.280 ;
        RECT 528.730 3.670 537.550 4.280 ;
        RECT 538.390 3.670 547.210 4.280 ;
        RECT 548.050 3.670 553.650 4.280 ;
        RECT 554.490 3.670 563.310 4.280 ;
        RECT 564.150 3.670 572.970 4.280 ;
        RECT 573.810 3.670 582.630 4.280 ;
        RECT 583.470 3.670 589.070 4.280 ;
        RECT 589.910 3.670 598.730 4.280 ;
        RECT 599.570 3.670 608.390 4.280 ;
        RECT 609.230 3.670 618.050 4.280 ;
        RECT 618.890 3.670 624.490 4.280 ;
        RECT 625.330 3.670 634.150 4.280 ;
        RECT 634.990 3.670 643.810 4.280 ;
        RECT 644.650 3.670 653.470 4.280 ;
        RECT 654.310 3.670 659.910 4.280 ;
        RECT 660.750 3.670 669.570 4.280 ;
        RECT 670.410 3.670 679.230 4.280 ;
        RECT 680.070 3.670 688.890 4.280 ;
        RECT 689.730 3.670 695.330 4.280 ;
        RECT 696.170 3.670 704.990 4.280 ;
        RECT 705.830 3.670 714.650 4.280 ;
        RECT 715.490 3.670 724.310 4.280 ;
        RECT 725.150 3.670 730.750 4.280 ;
        RECT 731.590 3.670 740.410 4.280 ;
        RECT 741.250 3.670 750.070 4.280 ;
        RECT 750.910 3.670 759.730 4.280 ;
        RECT 760.570 3.670 766.170 4.280 ;
        RECT 767.010 3.670 775.830 4.280 ;
        RECT 776.670 3.670 785.490 4.280 ;
        RECT 786.330 3.670 795.150 4.280 ;
        RECT 795.990 3.670 801.590 4.280 ;
        RECT 802.430 3.670 811.250 4.280 ;
        RECT 812.090 3.670 820.910 4.280 ;
        RECT 821.750 3.670 827.350 4.280 ;
        RECT 828.190 3.670 837.010 4.280 ;
        RECT 837.850 3.670 846.670 4.280 ;
        RECT 847.510 3.670 856.330 4.280 ;
        RECT 857.170 3.670 862.770 4.280 ;
        RECT 863.610 3.670 872.430 4.280 ;
        RECT 873.270 3.670 882.090 4.280 ;
        RECT 882.930 3.670 891.750 4.280 ;
        RECT 892.590 3.670 898.190 4.280 ;
        RECT 899.030 3.670 907.850 4.280 ;
        RECT 908.690 3.670 917.510 4.280 ;
        RECT 918.350 3.670 927.170 4.280 ;
        RECT 928.010 3.670 933.610 4.280 ;
        RECT 934.450 3.670 943.270 4.280 ;
        RECT 944.110 3.670 952.930 4.280 ;
        RECT 953.770 3.670 962.590 4.280 ;
        RECT 963.430 3.670 969.030 4.280 ;
        RECT 969.870 3.670 978.690 4.280 ;
        RECT 979.530 3.670 988.350 4.280 ;
        RECT 989.190 3.670 998.010 4.280 ;
        RECT 998.850 3.670 1004.450 4.280 ;
        RECT 1005.290 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1023.770 4.280 ;
        RECT 1024.610 3.670 1033.430 4.280 ;
        RECT 1034.270 3.670 1039.870 4.280 ;
        RECT 1040.710 3.670 1049.530 4.280 ;
        RECT 1050.370 3.670 1059.190 4.280 ;
        RECT 1060.030 3.670 1068.850 4.280 ;
        RECT 1069.690 3.670 1075.290 4.280 ;
        RECT 1076.130 3.670 1084.950 4.280 ;
        RECT 1085.790 3.670 1094.610 4.280 ;
        RECT 1095.450 3.670 1104.270 4.280 ;
        RECT 1105.110 3.670 1110.710 4.280 ;
        RECT 1111.550 3.670 1120.370 4.280 ;
        RECT 1121.210 3.670 1130.030 4.280 ;
        RECT 1130.870 3.670 1139.690 4.280 ;
        RECT 1140.530 3.670 1146.130 4.280 ;
        RECT 1146.970 3.670 1155.790 4.280 ;
        RECT 1156.630 3.670 1165.450 4.280 ;
        RECT 1166.290 3.670 1175.110 4.280 ;
        RECT 1175.950 3.670 1181.550 4.280 ;
        RECT 1182.390 3.670 1191.210 4.280 ;
        RECT 1192.050 3.670 1200.870 4.280 ;
        RECT 1201.710 3.670 1210.530 4.280 ;
        RECT 1211.370 3.670 1216.970 4.280 ;
        RECT 1217.810 3.670 1226.630 4.280 ;
        RECT 1227.470 3.670 1236.290 4.280 ;
        RECT 1237.130 3.670 1242.730 4.280 ;
        RECT 1243.570 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1262.050 4.280 ;
        RECT 1262.890 3.670 1271.710 4.280 ;
        RECT 1272.550 3.670 1278.150 4.280 ;
        RECT 1278.990 3.670 1287.810 4.280 ;
        RECT 1288.650 3.670 1297.470 4.280 ;
        RECT 1298.310 3.670 1307.130 4.280 ;
        RECT 1307.970 3.670 1313.570 4.280 ;
        RECT 1314.410 3.670 1323.230 4.280 ;
        RECT 1324.070 3.670 1332.890 4.280 ;
        RECT 1333.730 3.670 1342.550 4.280 ;
        RECT 1343.390 3.670 1348.990 4.280 ;
        RECT 1349.830 3.670 1358.650 4.280 ;
        RECT 1359.490 3.670 1368.310 4.280 ;
        RECT 1369.150 3.670 1377.970 4.280 ;
        RECT 1378.810 3.670 1384.410 4.280 ;
        RECT 1385.250 3.670 1394.070 4.280 ;
        RECT 1394.910 3.670 1403.730 4.280 ;
        RECT 1404.570 3.670 1413.390 4.280 ;
        RECT 1414.230 3.670 1419.830 4.280 ;
        RECT 1420.670 3.670 1429.490 4.280 ;
        RECT 1430.330 3.670 1439.150 4.280 ;
        RECT 1439.990 3.670 1448.810 4.280 ;
        RECT 1449.650 3.670 1455.250 4.280 ;
        RECT 1456.090 3.670 1464.910 4.280 ;
        RECT 1465.750 3.670 1474.570 4.280 ;
        RECT 1475.410 3.670 1484.230 4.280 ;
        RECT 1485.070 3.670 1490.670 4.280 ;
        RECT 1491.510 3.670 1500.330 4.280 ;
        RECT 1501.170 3.670 1509.990 4.280 ;
        RECT 1510.830 3.670 1519.650 4.280 ;
        RECT 1520.490 3.670 1526.090 4.280 ;
        RECT 1526.930 3.670 1535.750 4.280 ;
        RECT 1536.590 3.670 1545.410 4.280 ;
        RECT 1546.250 3.670 1555.070 4.280 ;
        RECT 1555.910 3.670 1561.510 4.280 ;
        RECT 1562.350 3.670 1571.170 4.280 ;
        RECT 1572.010 3.670 1580.830 4.280 ;
        RECT 1581.670 3.670 1590.130 4.280 ;
      LAYER met3 ;
        RECT 4.400 1135.240 1595.600 1136.105 ;
        RECT 4.000 1129.840 1596.000 1135.240 ;
        RECT 4.400 1128.440 1596.000 1129.840 ;
        RECT 4.000 1126.440 1596.000 1128.440 ;
        RECT 4.000 1125.040 1595.600 1126.440 ;
        RECT 4.000 1119.640 1596.000 1125.040 ;
        RECT 4.400 1118.240 1595.600 1119.640 ;
        RECT 4.000 1109.440 1596.000 1118.240 ;
        RECT 4.400 1108.040 1595.600 1109.440 ;
        RECT 4.000 1099.240 1596.000 1108.040 ;
        RECT 4.400 1097.840 1595.600 1099.240 ;
        RECT 4.000 1092.440 1596.000 1097.840 ;
        RECT 4.400 1091.040 1596.000 1092.440 ;
        RECT 4.000 1089.040 1596.000 1091.040 ;
        RECT 4.000 1087.640 1595.600 1089.040 ;
        RECT 4.000 1082.240 1596.000 1087.640 ;
        RECT 4.400 1080.840 1595.600 1082.240 ;
        RECT 4.000 1072.040 1596.000 1080.840 ;
        RECT 4.400 1070.640 1595.600 1072.040 ;
        RECT 4.000 1061.840 1596.000 1070.640 ;
        RECT 4.400 1060.440 1595.600 1061.840 ;
        RECT 4.000 1055.040 1596.000 1060.440 ;
        RECT 4.400 1053.640 1596.000 1055.040 ;
        RECT 4.000 1051.640 1596.000 1053.640 ;
        RECT 4.000 1050.240 1595.600 1051.640 ;
        RECT 4.000 1044.840 1596.000 1050.240 ;
        RECT 4.400 1043.440 1595.600 1044.840 ;
        RECT 4.000 1034.640 1596.000 1043.440 ;
        RECT 4.400 1033.240 1595.600 1034.640 ;
        RECT 4.000 1024.440 1596.000 1033.240 ;
        RECT 4.400 1023.040 1595.600 1024.440 ;
        RECT 4.000 1017.640 1596.000 1023.040 ;
        RECT 4.400 1016.240 1596.000 1017.640 ;
        RECT 4.000 1014.240 1596.000 1016.240 ;
        RECT 4.000 1012.840 1595.600 1014.240 ;
        RECT 4.000 1007.440 1596.000 1012.840 ;
        RECT 4.400 1006.040 1595.600 1007.440 ;
        RECT 4.000 997.240 1596.000 1006.040 ;
        RECT 4.400 995.840 1595.600 997.240 ;
        RECT 4.000 987.040 1596.000 995.840 ;
        RECT 4.400 985.640 1595.600 987.040 ;
        RECT 4.000 980.240 1596.000 985.640 ;
        RECT 4.400 978.840 1596.000 980.240 ;
        RECT 4.000 976.840 1596.000 978.840 ;
        RECT 4.000 975.440 1595.600 976.840 ;
        RECT 4.000 970.040 1596.000 975.440 ;
        RECT 4.400 968.640 1595.600 970.040 ;
        RECT 4.000 959.840 1596.000 968.640 ;
        RECT 4.400 958.440 1595.600 959.840 ;
        RECT 4.000 949.640 1596.000 958.440 ;
        RECT 4.400 948.240 1595.600 949.640 ;
        RECT 4.000 942.840 1596.000 948.240 ;
        RECT 4.400 941.440 1596.000 942.840 ;
        RECT 4.000 939.440 1596.000 941.440 ;
        RECT 4.000 938.040 1595.600 939.440 ;
        RECT 4.000 932.640 1596.000 938.040 ;
        RECT 4.400 931.240 1595.600 932.640 ;
        RECT 4.000 922.440 1596.000 931.240 ;
        RECT 4.400 921.040 1595.600 922.440 ;
        RECT 4.000 912.240 1596.000 921.040 ;
        RECT 4.400 910.840 1595.600 912.240 ;
        RECT 4.000 905.440 1596.000 910.840 ;
        RECT 4.400 904.040 1595.600 905.440 ;
        RECT 4.000 895.240 1596.000 904.040 ;
        RECT 4.400 893.840 1595.600 895.240 ;
        RECT 4.000 885.040 1596.000 893.840 ;
        RECT 4.400 883.640 1595.600 885.040 ;
        RECT 4.000 874.840 1596.000 883.640 ;
        RECT 4.400 873.440 1595.600 874.840 ;
        RECT 4.000 868.040 1596.000 873.440 ;
        RECT 4.400 866.640 1595.600 868.040 ;
        RECT 4.000 857.840 1596.000 866.640 ;
        RECT 4.400 856.440 1595.600 857.840 ;
        RECT 4.000 847.640 1596.000 856.440 ;
        RECT 4.400 846.240 1595.600 847.640 ;
        RECT 4.000 840.840 1596.000 846.240 ;
        RECT 4.400 839.440 1596.000 840.840 ;
        RECT 4.000 837.440 1596.000 839.440 ;
        RECT 4.000 836.040 1595.600 837.440 ;
        RECT 4.000 830.640 1596.000 836.040 ;
        RECT 4.400 829.240 1595.600 830.640 ;
        RECT 4.000 820.440 1596.000 829.240 ;
        RECT 4.400 819.040 1595.600 820.440 ;
        RECT 4.000 810.240 1596.000 819.040 ;
        RECT 4.400 808.840 1595.600 810.240 ;
        RECT 4.000 803.440 1596.000 808.840 ;
        RECT 4.400 802.040 1596.000 803.440 ;
        RECT 4.000 800.040 1596.000 802.040 ;
        RECT 4.000 798.640 1595.600 800.040 ;
        RECT 4.000 793.240 1596.000 798.640 ;
        RECT 4.400 791.840 1595.600 793.240 ;
        RECT 4.000 783.040 1596.000 791.840 ;
        RECT 4.400 781.640 1595.600 783.040 ;
        RECT 4.000 772.840 1596.000 781.640 ;
        RECT 4.400 771.440 1595.600 772.840 ;
        RECT 4.000 766.040 1596.000 771.440 ;
        RECT 4.400 764.640 1596.000 766.040 ;
        RECT 4.000 762.640 1596.000 764.640 ;
        RECT 4.000 761.240 1595.600 762.640 ;
        RECT 4.000 755.840 1596.000 761.240 ;
        RECT 4.400 754.440 1595.600 755.840 ;
        RECT 4.000 745.640 1596.000 754.440 ;
        RECT 4.400 744.240 1595.600 745.640 ;
        RECT 4.000 735.440 1596.000 744.240 ;
        RECT 4.400 734.040 1595.600 735.440 ;
        RECT 4.000 728.640 1596.000 734.040 ;
        RECT 4.400 727.240 1596.000 728.640 ;
        RECT 4.000 725.240 1596.000 727.240 ;
        RECT 4.000 723.840 1595.600 725.240 ;
        RECT 4.000 718.440 1596.000 723.840 ;
        RECT 4.400 717.040 1595.600 718.440 ;
        RECT 4.000 708.240 1596.000 717.040 ;
        RECT 4.400 706.840 1595.600 708.240 ;
        RECT 4.000 698.040 1596.000 706.840 ;
        RECT 4.400 696.640 1595.600 698.040 ;
        RECT 4.000 691.240 1596.000 696.640 ;
        RECT 4.400 689.840 1596.000 691.240 ;
        RECT 4.000 687.840 1596.000 689.840 ;
        RECT 4.000 686.440 1595.600 687.840 ;
        RECT 4.000 681.040 1596.000 686.440 ;
        RECT 4.400 679.640 1595.600 681.040 ;
        RECT 4.000 670.840 1596.000 679.640 ;
        RECT 4.400 669.440 1595.600 670.840 ;
        RECT 4.000 660.640 1596.000 669.440 ;
        RECT 4.400 659.240 1595.600 660.640 ;
        RECT 4.000 653.840 1596.000 659.240 ;
        RECT 4.400 652.440 1596.000 653.840 ;
        RECT 4.000 650.440 1596.000 652.440 ;
        RECT 4.000 649.040 1595.600 650.440 ;
        RECT 4.000 643.640 1596.000 649.040 ;
        RECT 4.400 642.240 1595.600 643.640 ;
        RECT 4.000 633.440 1596.000 642.240 ;
        RECT 4.400 632.040 1595.600 633.440 ;
        RECT 4.000 623.240 1596.000 632.040 ;
        RECT 4.400 621.840 1595.600 623.240 ;
        RECT 4.000 616.440 1596.000 621.840 ;
        RECT 4.400 615.040 1596.000 616.440 ;
        RECT 4.000 613.040 1596.000 615.040 ;
        RECT 4.000 611.640 1595.600 613.040 ;
        RECT 4.000 606.240 1596.000 611.640 ;
        RECT 4.400 604.840 1595.600 606.240 ;
        RECT 4.000 596.040 1596.000 604.840 ;
        RECT 4.400 594.640 1595.600 596.040 ;
        RECT 4.000 585.840 1596.000 594.640 ;
        RECT 4.400 584.440 1595.600 585.840 ;
        RECT 4.000 579.040 1596.000 584.440 ;
        RECT 4.400 577.640 1596.000 579.040 ;
        RECT 4.000 575.640 1596.000 577.640 ;
        RECT 4.000 574.240 1595.600 575.640 ;
        RECT 4.000 568.840 1596.000 574.240 ;
        RECT 4.400 567.440 1595.600 568.840 ;
        RECT 4.000 558.640 1596.000 567.440 ;
        RECT 4.400 557.240 1595.600 558.640 ;
        RECT 4.000 548.440 1596.000 557.240 ;
        RECT 4.400 547.040 1595.600 548.440 ;
        RECT 4.000 541.640 1596.000 547.040 ;
        RECT 4.400 540.240 1596.000 541.640 ;
        RECT 4.000 538.240 1596.000 540.240 ;
        RECT 4.000 536.840 1595.600 538.240 ;
        RECT 4.000 531.440 1596.000 536.840 ;
        RECT 4.400 530.040 1595.600 531.440 ;
        RECT 4.000 521.240 1596.000 530.040 ;
        RECT 4.400 519.840 1595.600 521.240 ;
        RECT 4.000 511.040 1596.000 519.840 ;
        RECT 4.400 509.640 1595.600 511.040 ;
        RECT 4.000 504.240 1596.000 509.640 ;
        RECT 4.400 502.840 1596.000 504.240 ;
        RECT 4.000 500.840 1596.000 502.840 ;
        RECT 4.000 499.440 1595.600 500.840 ;
        RECT 4.000 494.040 1596.000 499.440 ;
        RECT 4.400 492.640 1595.600 494.040 ;
        RECT 4.000 483.840 1596.000 492.640 ;
        RECT 4.400 482.440 1595.600 483.840 ;
        RECT 4.000 473.640 1596.000 482.440 ;
        RECT 4.400 472.240 1595.600 473.640 ;
        RECT 4.000 466.840 1596.000 472.240 ;
        RECT 4.400 465.440 1595.600 466.840 ;
        RECT 4.000 456.640 1596.000 465.440 ;
        RECT 4.400 455.240 1595.600 456.640 ;
        RECT 4.000 446.440 1596.000 455.240 ;
        RECT 4.400 445.040 1595.600 446.440 ;
        RECT 4.000 436.240 1596.000 445.040 ;
        RECT 4.400 434.840 1595.600 436.240 ;
        RECT 4.000 429.440 1596.000 434.840 ;
        RECT 4.400 428.040 1595.600 429.440 ;
        RECT 4.000 419.240 1596.000 428.040 ;
        RECT 4.400 417.840 1595.600 419.240 ;
        RECT 4.000 409.040 1596.000 417.840 ;
        RECT 4.400 407.640 1595.600 409.040 ;
        RECT 4.000 402.240 1596.000 407.640 ;
        RECT 4.400 400.840 1596.000 402.240 ;
        RECT 4.000 398.840 1596.000 400.840 ;
        RECT 4.000 397.440 1595.600 398.840 ;
        RECT 4.000 392.040 1596.000 397.440 ;
        RECT 4.400 390.640 1595.600 392.040 ;
        RECT 4.000 381.840 1596.000 390.640 ;
        RECT 4.400 380.440 1595.600 381.840 ;
        RECT 4.000 371.640 1596.000 380.440 ;
        RECT 4.400 370.240 1595.600 371.640 ;
        RECT 4.000 364.840 1596.000 370.240 ;
        RECT 4.400 363.440 1596.000 364.840 ;
        RECT 4.000 361.440 1596.000 363.440 ;
        RECT 4.000 360.040 1595.600 361.440 ;
        RECT 4.000 354.640 1596.000 360.040 ;
        RECT 4.400 353.240 1595.600 354.640 ;
        RECT 4.000 344.440 1596.000 353.240 ;
        RECT 4.400 343.040 1595.600 344.440 ;
        RECT 4.000 334.240 1596.000 343.040 ;
        RECT 4.400 332.840 1595.600 334.240 ;
        RECT 4.000 327.440 1596.000 332.840 ;
        RECT 4.400 326.040 1596.000 327.440 ;
        RECT 4.000 324.040 1596.000 326.040 ;
        RECT 4.000 322.640 1595.600 324.040 ;
        RECT 4.000 317.240 1596.000 322.640 ;
        RECT 4.400 315.840 1595.600 317.240 ;
        RECT 4.000 307.040 1596.000 315.840 ;
        RECT 4.400 305.640 1595.600 307.040 ;
        RECT 4.000 296.840 1596.000 305.640 ;
        RECT 4.400 295.440 1595.600 296.840 ;
        RECT 4.000 290.040 1596.000 295.440 ;
        RECT 4.400 288.640 1596.000 290.040 ;
        RECT 4.000 286.640 1596.000 288.640 ;
        RECT 4.000 285.240 1595.600 286.640 ;
        RECT 4.000 279.840 1596.000 285.240 ;
        RECT 4.400 278.440 1595.600 279.840 ;
        RECT 4.000 269.640 1596.000 278.440 ;
        RECT 4.400 268.240 1595.600 269.640 ;
        RECT 4.000 259.440 1596.000 268.240 ;
        RECT 4.400 258.040 1595.600 259.440 ;
        RECT 4.000 252.640 1596.000 258.040 ;
        RECT 4.400 251.240 1596.000 252.640 ;
        RECT 4.000 249.240 1596.000 251.240 ;
        RECT 4.000 247.840 1595.600 249.240 ;
        RECT 4.000 242.440 1596.000 247.840 ;
        RECT 4.400 241.040 1595.600 242.440 ;
        RECT 4.000 232.240 1596.000 241.040 ;
        RECT 4.400 230.840 1595.600 232.240 ;
        RECT 4.000 222.040 1596.000 230.840 ;
        RECT 4.400 220.640 1595.600 222.040 ;
        RECT 4.000 215.240 1596.000 220.640 ;
        RECT 4.400 213.840 1596.000 215.240 ;
        RECT 4.000 211.840 1596.000 213.840 ;
        RECT 4.000 210.440 1595.600 211.840 ;
        RECT 4.000 205.040 1596.000 210.440 ;
        RECT 4.400 203.640 1595.600 205.040 ;
        RECT 4.000 194.840 1596.000 203.640 ;
        RECT 4.400 193.440 1595.600 194.840 ;
        RECT 4.000 184.640 1596.000 193.440 ;
        RECT 4.400 183.240 1595.600 184.640 ;
        RECT 4.000 177.840 1596.000 183.240 ;
        RECT 4.400 176.440 1596.000 177.840 ;
        RECT 4.000 174.440 1596.000 176.440 ;
        RECT 4.000 173.040 1595.600 174.440 ;
        RECT 4.000 167.640 1596.000 173.040 ;
        RECT 4.400 166.240 1595.600 167.640 ;
        RECT 4.000 157.440 1596.000 166.240 ;
        RECT 4.400 156.040 1595.600 157.440 ;
        RECT 4.000 147.240 1596.000 156.040 ;
        RECT 4.400 145.840 1595.600 147.240 ;
        RECT 4.000 140.440 1596.000 145.840 ;
        RECT 4.400 139.040 1596.000 140.440 ;
        RECT 4.000 137.040 1596.000 139.040 ;
        RECT 4.000 135.640 1595.600 137.040 ;
        RECT 4.000 130.240 1596.000 135.640 ;
        RECT 4.400 128.840 1595.600 130.240 ;
        RECT 4.000 120.040 1596.000 128.840 ;
        RECT 4.400 118.640 1595.600 120.040 ;
        RECT 4.000 109.840 1596.000 118.640 ;
        RECT 4.400 108.440 1595.600 109.840 ;
        RECT 4.000 103.040 1596.000 108.440 ;
        RECT 4.400 101.640 1596.000 103.040 ;
        RECT 4.000 99.640 1596.000 101.640 ;
        RECT 4.000 98.240 1595.600 99.640 ;
        RECT 4.000 92.840 1596.000 98.240 ;
        RECT 4.400 91.440 1595.600 92.840 ;
        RECT 4.000 82.640 1596.000 91.440 ;
        RECT 4.400 81.240 1595.600 82.640 ;
        RECT 4.000 72.440 1596.000 81.240 ;
        RECT 4.400 71.040 1595.600 72.440 ;
        RECT 4.000 65.640 1596.000 71.040 ;
        RECT 4.400 64.240 1596.000 65.640 ;
        RECT 4.000 62.240 1596.000 64.240 ;
        RECT 4.000 60.840 1595.600 62.240 ;
        RECT 4.000 55.440 1596.000 60.840 ;
        RECT 4.400 54.040 1595.600 55.440 ;
        RECT 4.000 45.240 1596.000 54.040 ;
        RECT 4.400 43.840 1595.600 45.240 ;
        RECT 4.000 35.040 1596.000 43.840 ;
        RECT 4.400 33.640 1595.600 35.040 ;
        RECT 4.000 28.240 1596.000 33.640 ;
        RECT 4.400 26.840 1595.600 28.240 ;
        RECT 4.000 18.040 1596.000 26.840 ;
        RECT 4.400 16.640 1595.600 18.040 ;
        RECT 4.000 10.715 1596.000 16.640 ;
      LAYER met4 ;
        RECT 194.415 1026.860 220.640 1035.465 ;
        RECT 223.040 1026.860 270.640 1035.465 ;
        RECT 273.040 1026.860 320.640 1035.465 ;
        RECT 323.040 1026.860 370.640 1035.465 ;
        RECT 373.040 1026.860 420.640 1035.465 ;
        RECT 423.040 1026.860 470.640 1035.465 ;
        RECT 473.040 1026.860 520.640 1035.465 ;
        RECT 523.040 1026.860 570.640 1035.465 ;
        RECT 573.040 1026.860 620.640 1035.465 ;
        RECT 623.040 1026.860 670.640 1035.465 ;
        RECT 673.040 1026.860 720.640 1035.465 ;
        RECT 194.415 610.640 720.640 1026.860 ;
        RECT 194.415 506.860 220.640 610.640 ;
        RECT 223.040 506.860 270.640 610.640 ;
        RECT 273.040 506.860 320.640 610.640 ;
        RECT 323.040 506.860 370.640 610.640 ;
        RECT 373.040 506.860 420.640 610.640 ;
        RECT 423.040 506.860 470.640 610.640 ;
        RECT 473.040 506.860 520.640 610.640 ;
        RECT 523.040 506.860 570.640 610.640 ;
        RECT 573.040 506.860 620.640 610.640 ;
        RECT 623.040 506.860 670.640 610.640 ;
        RECT 673.040 506.860 720.640 610.640 ;
        RECT 194.415 90.640 720.640 506.860 ;
        RECT 194.415 83.135 220.640 90.640 ;
        RECT 223.040 83.135 270.640 90.640 ;
        RECT 273.040 83.135 320.640 90.640 ;
        RECT 323.040 83.135 370.640 90.640 ;
        RECT 373.040 83.135 420.640 90.640 ;
        RECT 423.040 83.135 470.640 90.640 ;
        RECT 473.040 83.135 520.640 90.640 ;
        RECT 523.040 83.135 570.640 90.640 ;
        RECT 573.040 83.135 620.640 90.640 ;
        RECT 623.040 83.135 670.640 90.640 ;
        RECT 673.040 83.135 720.640 90.640 ;
        RECT 723.040 83.135 770.640 1035.465 ;
        RECT 773.040 83.135 820.640 1035.465 ;
        RECT 823.040 83.135 870.640 1035.465 ;
        RECT 873.040 1026.860 920.640 1035.465 ;
        RECT 923.040 1026.860 970.640 1035.465 ;
        RECT 973.040 1026.860 1020.640 1035.465 ;
        RECT 1023.040 1026.860 1070.640 1035.465 ;
        RECT 1073.040 1026.860 1120.640 1035.465 ;
        RECT 1123.040 1026.860 1170.640 1035.465 ;
        RECT 1173.040 1026.860 1220.640 1035.465 ;
        RECT 1223.040 1026.860 1270.640 1035.465 ;
        RECT 1273.040 1026.860 1320.640 1035.465 ;
        RECT 1323.040 1026.860 1370.640 1035.465 ;
        RECT 1373.040 1026.860 1383.385 1035.465 ;
        RECT 873.040 610.640 1383.385 1026.860 ;
        RECT 873.040 506.860 920.640 610.640 ;
        RECT 923.040 506.860 970.640 610.640 ;
        RECT 973.040 506.860 1020.640 610.640 ;
        RECT 1023.040 506.860 1070.640 610.640 ;
        RECT 1073.040 506.860 1120.640 610.640 ;
        RECT 1123.040 506.860 1170.640 610.640 ;
        RECT 1173.040 506.860 1220.640 610.640 ;
        RECT 1223.040 506.860 1270.640 610.640 ;
        RECT 1273.040 506.860 1320.640 610.640 ;
        RECT 1323.040 506.860 1370.640 610.640 ;
        RECT 1373.040 506.860 1383.385 610.640 ;
        RECT 873.040 90.640 1383.385 506.860 ;
        RECT 873.040 83.135 920.640 90.640 ;
        RECT 923.040 83.135 970.640 90.640 ;
        RECT 973.040 83.135 1020.640 90.640 ;
        RECT 1023.040 83.135 1070.640 90.640 ;
        RECT 1073.040 83.135 1120.640 90.640 ;
        RECT 1123.040 83.135 1170.640 90.640 ;
        RECT 1173.040 83.135 1220.640 90.640 ;
        RECT 1223.040 83.135 1270.640 90.640 ;
        RECT 1273.040 83.135 1320.640 90.640 ;
        RECT 1323.040 83.135 1370.640 90.640 ;
        RECT 1373.040 83.135 1383.385 90.640 ;
  END
END openram_demo
END LIBRARY

