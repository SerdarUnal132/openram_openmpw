magic
tech sky130A
magscale 1 2
timestamp 1653355972
<< obsli1 >>
rect 1104 2159 318872 225777
<< obsm1 >>
rect 14 2128 318872 225808
<< metal2 >>
rect 662 227200 718 228000
rect 2594 227200 2650 228000
rect 4526 227200 4582 228000
rect 5814 227200 5870 228000
rect 7746 227200 7802 228000
rect 9678 227200 9734 228000
rect 11610 227200 11666 228000
rect 12898 227200 12954 228000
rect 14830 227200 14886 228000
rect 16762 227200 16818 228000
rect 18694 227200 18750 228000
rect 19982 227200 20038 228000
rect 21914 227200 21970 228000
rect 23846 227200 23902 228000
rect 25778 227200 25834 228000
rect 27066 227200 27122 228000
rect 28998 227200 29054 228000
rect 30930 227200 30986 228000
rect 32218 227200 32274 228000
rect 34150 227200 34206 228000
rect 36082 227200 36138 228000
rect 38014 227200 38070 228000
rect 39302 227200 39358 228000
rect 41234 227200 41290 228000
rect 43166 227200 43222 228000
rect 45098 227200 45154 228000
rect 46386 227200 46442 228000
rect 48318 227200 48374 228000
rect 50250 227200 50306 228000
rect 52182 227200 52238 228000
rect 53470 227200 53526 228000
rect 55402 227200 55458 228000
rect 57334 227200 57390 228000
rect 59266 227200 59322 228000
rect 60554 227200 60610 228000
rect 62486 227200 62542 228000
rect 64418 227200 64474 228000
rect 66350 227200 66406 228000
rect 67638 227200 67694 228000
rect 69570 227200 69626 228000
rect 71502 227200 71558 228000
rect 73434 227200 73490 228000
rect 74722 227200 74778 228000
rect 76654 227200 76710 228000
rect 78586 227200 78642 228000
rect 80518 227200 80574 228000
rect 81806 227200 81862 228000
rect 83738 227200 83794 228000
rect 85670 227200 85726 228000
rect 87602 227200 87658 228000
rect 88890 227200 88946 228000
rect 90822 227200 90878 228000
rect 92754 227200 92810 228000
rect 94686 227200 94742 228000
rect 95974 227200 96030 228000
rect 97906 227200 97962 228000
rect 99838 227200 99894 228000
rect 101770 227200 101826 228000
rect 103058 227200 103114 228000
rect 104990 227200 105046 228000
rect 106922 227200 106978 228000
rect 108854 227200 108910 228000
rect 110142 227200 110198 228000
rect 112074 227200 112130 228000
rect 114006 227200 114062 228000
rect 115294 227200 115350 228000
rect 117226 227200 117282 228000
rect 119158 227200 119214 228000
rect 121090 227200 121146 228000
rect 122378 227200 122434 228000
rect 124310 227200 124366 228000
rect 126242 227200 126298 228000
rect 128174 227200 128230 228000
rect 129462 227200 129518 228000
rect 131394 227200 131450 228000
rect 133326 227200 133382 228000
rect 135258 227200 135314 228000
rect 136546 227200 136602 228000
rect 138478 227200 138534 228000
rect 140410 227200 140466 228000
rect 142342 227200 142398 228000
rect 143630 227200 143686 228000
rect 145562 227200 145618 228000
rect 147494 227200 147550 228000
rect 149426 227200 149482 228000
rect 150714 227200 150770 228000
rect 152646 227200 152702 228000
rect 154578 227200 154634 228000
rect 156510 227200 156566 228000
rect 157798 227200 157854 228000
rect 159730 227200 159786 228000
rect 161662 227200 161718 228000
rect 163594 227200 163650 228000
rect 164882 227200 164938 228000
rect 166814 227200 166870 228000
rect 168746 227200 168802 228000
rect 170678 227200 170734 228000
rect 171966 227200 172022 228000
rect 173898 227200 173954 228000
rect 175830 227200 175886 228000
rect 177762 227200 177818 228000
rect 179050 227200 179106 228000
rect 180982 227200 181038 228000
rect 182914 227200 182970 228000
rect 184846 227200 184902 228000
rect 186134 227200 186190 228000
rect 188066 227200 188122 228000
rect 189998 227200 190054 228000
rect 191930 227200 191986 228000
rect 193218 227200 193274 228000
rect 195150 227200 195206 228000
rect 197082 227200 197138 228000
rect 198370 227200 198426 228000
rect 200302 227200 200358 228000
rect 202234 227200 202290 228000
rect 204166 227200 204222 228000
rect 205454 227200 205510 228000
rect 207386 227200 207442 228000
rect 209318 227200 209374 228000
rect 211250 227200 211306 228000
rect 212538 227200 212594 228000
rect 214470 227200 214526 228000
rect 216402 227200 216458 228000
rect 218334 227200 218390 228000
rect 219622 227200 219678 228000
rect 221554 227200 221610 228000
rect 223486 227200 223542 228000
rect 225418 227200 225474 228000
rect 226706 227200 226762 228000
rect 228638 227200 228694 228000
rect 230570 227200 230626 228000
rect 232502 227200 232558 228000
rect 233790 227200 233846 228000
rect 235722 227200 235778 228000
rect 237654 227200 237710 228000
rect 239586 227200 239642 228000
rect 240874 227200 240930 228000
rect 242806 227200 242862 228000
rect 244738 227200 244794 228000
rect 246670 227200 246726 228000
rect 247958 227200 248014 228000
rect 249890 227200 249946 228000
rect 251822 227200 251878 228000
rect 253754 227200 253810 228000
rect 255042 227200 255098 228000
rect 256974 227200 257030 228000
rect 258906 227200 258962 228000
rect 260838 227200 260894 228000
rect 262126 227200 262182 228000
rect 264058 227200 264114 228000
rect 265990 227200 266046 228000
rect 267922 227200 267978 228000
rect 269210 227200 269266 228000
rect 271142 227200 271198 228000
rect 273074 227200 273130 228000
rect 275006 227200 275062 228000
rect 276294 227200 276350 228000
rect 278226 227200 278282 228000
rect 280158 227200 280214 228000
rect 281446 227200 281502 228000
rect 283378 227200 283434 228000
rect 285310 227200 285366 228000
rect 287242 227200 287298 228000
rect 288530 227200 288586 228000
rect 290462 227200 290518 228000
rect 292394 227200 292450 228000
rect 294326 227200 294382 228000
rect 295614 227200 295670 228000
rect 297546 227200 297602 228000
rect 299478 227200 299534 228000
rect 301410 227200 301466 228000
rect 302698 227200 302754 228000
rect 304630 227200 304686 228000
rect 306562 227200 306618 228000
rect 308494 227200 308550 228000
rect 309782 227200 309838 228000
rect 311714 227200 311770 228000
rect 313646 227200 313702 228000
rect 315578 227200 315634 228000
rect 316866 227200 316922 228000
rect 318798 227200 318854 228000
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36726 0 36782 800
rect 38658 0 38714 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 50894 0 50950 800
rect 52826 0 52882 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 59910 0 59966 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 65062 0 65118 800
rect 66994 0 67050 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 72146 0 72202 800
rect 74078 0 74134 800
rect 76010 0 76066 800
rect 77298 0 77354 800
rect 79230 0 79286 800
rect 81162 0 81218 800
rect 82450 0 82506 800
rect 84382 0 84438 800
rect 86314 0 86370 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 91466 0 91522 800
rect 93398 0 93454 800
rect 95330 0 95386 800
rect 96618 0 96674 800
rect 98550 0 98606 800
rect 100482 0 100538 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 105634 0 105690 800
rect 107566 0 107622 800
rect 109498 0 109554 800
rect 110786 0 110842 800
rect 112718 0 112774 800
rect 114650 0 114706 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 119802 0 119858 800
rect 121734 0 121790 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 126886 0 126942 800
rect 128818 0 128874 800
rect 130750 0 130806 800
rect 132038 0 132094 800
rect 133970 0 134026 800
rect 135902 0 135958 800
rect 137834 0 137890 800
rect 139122 0 139178 800
rect 141054 0 141110 800
rect 142986 0 143042 800
rect 144918 0 144974 800
rect 146206 0 146262 800
rect 148138 0 148194 800
rect 150070 0 150126 800
rect 152002 0 152058 800
rect 153290 0 153346 800
rect 155222 0 155278 800
rect 157154 0 157210 800
rect 159086 0 159142 800
rect 160374 0 160430 800
rect 162306 0 162362 800
rect 164238 0 164294 800
rect 165526 0 165582 800
rect 167458 0 167514 800
rect 169390 0 169446 800
rect 171322 0 171378 800
rect 172610 0 172666 800
rect 174542 0 174598 800
rect 176474 0 176530 800
rect 178406 0 178462 800
rect 179694 0 179750 800
rect 181626 0 181682 800
rect 183558 0 183614 800
rect 185490 0 185546 800
rect 186778 0 186834 800
rect 188710 0 188766 800
rect 190642 0 190698 800
rect 192574 0 192630 800
rect 193862 0 193918 800
rect 195794 0 195850 800
rect 197726 0 197782 800
rect 199658 0 199714 800
rect 200946 0 201002 800
rect 202878 0 202934 800
rect 204810 0 204866 800
rect 206742 0 206798 800
rect 208030 0 208086 800
rect 209962 0 210018 800
rect 211894 0 211950 800
rect 213826 0 213882 800
rect 215114 0 215170 800
rect 217046 0 217102 800
rect 218978 0 219034 800
rect 220910 0 220966 800
rect 222198 0 222254 800
rect 224130 0 224186 800
rect 226062 0 226118 800
rect 227994 0 228050 800
rect 229282 0 229338 800
rect 231214 0 231270 800
rect 233146 0 233202 800
rect 235078 0 235134 800
rect 236366 0 236422 800
rect 238298 0 238354 800
rect 240230 0 240286 800
rect 242162 0 242218 800
rect 243450 0 243506 800
rect 245382 0 245438 800
rect 247314 0 247370 800
rect 248602 0 248658 800
rect 250534 0 250590 800
rect 252466 0 252522 800
rect 254398 0 254454 800
rect 255686 0 255742 800
rect 257618 0 257674 800
rect 259550 0 259606 800
rect 261482 0 261538 800
rect 262770 0 262826 800
rect 264702 0 264758 800
rect 266634 0 266690 800
rect 268566 0 268622 800
rect 269854 0 269910 800
rect 271786 0 271842 800
rect 273718 0 273774 800
rect 275650 0 275706 800
rect 276938 0 276994 800
rect 278870 0 278926 800
rect 280802 0 280858 800
rect 282734 0 282790 800
rect 284022 0 284078 800
rect 285954 0 286010 800
rect 287886 0 287942 800
rect 289818 0 289874 800
rect 291106 0 291162 800
rect 293038 0 293094 800
rect 294970 0 295026 800
rect 296902 0 296958 800
rect 298190 0 298246 800
rect 300122 0 300178 800
rect 302054 0 302110 800
rect 303986 0 304042 800
rect 305274 0 305330 800
rect 307206 0 307262 800
rect 309138 0 309194 800
rect 311070 0 311126 800
rect 312358 0 312414 800
rect 314290 0 314346 800
rect 316222 0 316278 800
rect 318154 0 318210 800
rect 319442 0 319498 800
<< obsm2 >>
rect 20 227144 606 227338
rect 774 227144 2538 227338
rect 2706 227144 4470 227338
rect 4638 227144 5758 227338
rect 5926 227144 7690 227338
rect 7858 227144 9622 227338
rect 9790 227144 11554 227338
rect 11722 227144 12842 227338
rect 13010 227144 14774 227338
rect 14942 227144 16706 227338
rect 16874 227144 18638 227338
rect 18806 227144 19926 227338
rect 20094 227144 21858 227338
rect 22026 227144 23790 227338
rect 23958 227144 25722 227338
rect 25890 227144 27010 227338
rect 27178 227144 28942 227338
rect 29110 227144 30874 227338
rect 31042 227144 32162 227338
rect 32330 227144 34094 227338
rect 34262 227144 36026 227338
rect 36194 227144 37958 227338
rect 38126 227144 39246 227338
rect 39414 227144 41178 227338
rect 41346 227144 43110 227338
rect 43278 227144 45042 227338
rect 45210 227144 46330 227338
rect 46498 227144 48262 227338
rect 48430 227144 50194 227338
rect 50362 227144 52126 227338
rect 52294 227144 53414 227338
rect 53582 227144 55346 227338
rect 55514 227144 57278 227338
rect 57446 227144 59210 227338
rect 59378 227144 60498 227338
rect 60666 227144 62430 227338
rect 62598 227144 64362 227338
rect 64530 227144 66294 227338
rect 66462 227144 67582 227338
rect 67750 227144 69514 227338
rect 69682 227144 71446 227338
rect 71614 227144 73378 227338
rect 73546 227144 74666 227338
rect 74834 227144 76598 227338
rect 76766 227144 78530 227338
rect 78698 227144 80462 227338
rect 80630 227144 81750 227338
rect 81918 227144 83682 227338
rect 83850 227144 85614 227338
rect 85782 227144 87546 227338
rect 87714 227144 88834 227338
rect 89002 227144 90766 227338
rect 90934 227144 92698 227338
rect 92866 227144 94630 227338
rect 94798 227144 95918 227338
rect 96086 227144 97850 227338
rect 98018 227144 99782 227338
rect 99950 227144 101714 227338
rect 101882 227144 103002 227338
rect 103170 227144 104934 227338
rect 105102 227144 106866 227338
rect 107034 227144 108798 227338
rect 108966 227144 110086 227338
rect 110254 227144 112018 227338
rect 112186 227144 113950 227338
rect 114118 227144 115238 227338
rect 115406 227144 117170 227338
rect 117338 227144 119102 227338
rect 119270 227144 121034 227338
rect 121202 227144 122322 227338
rect 122490 227144 124254 227338
rect 124422 227144 126186 227338
rect 126354 227144 128118 227338
rect 128286 227144 129406 227338
rect 129574 227144 131338 227338
rect 131506 227144 133270 227338
rect 133438 227144 135202 227338
rect 135370 227144 136490 227338
rect 136658 227144 138422 227338
rect 138590 227144 140354 227338
rect 140522 227144 142286 227338
rect 142454 227144 143574 227338
rect 143742 227144 145506 227338
rect 145674 227144 147438 227338
rect 147606 227144 149370 227338
rect 149538 227144 150658 227338
rect 150826 227144 152590 227338
rect 152758 227144 154522 227338
rect 154690 227144 156454 227338
rect 156622 227144 157742 227338
rect 157910 227144 159674 227338
rect 159842 227144 161606 227338
rect 161774 227144 163538 227338
rect 163706 227144 164826 227338
rect 164994 227144 166758 227338
rect 166926 227144 168690 227338
rect 168858 227144 170622 227338
rect 170790 227144 171910 227338
rect 172078 227144 173842 227338
rect 174010 227144 175774 227338
rect 175942 227144 177706 227338
rect 177874 227144 178994 227338
rect 179162 227144 180926 227338
rect 181094 227144 182858 227338
rect 183026 227144 184790 227338
rect 184958 227144 186078 227338
rect 186246 227144 188010 227338
rect 188178 227144 189942 227338
rect 190110 227144 191874 227338
rect 192042 227144 193162 227338
rect 193330 227144 195094 227338
rect 195262 227144 197026 227338
rect 197194 227144 198314 227338
rect 198482 227144 200246 227338
rect 200414 227144 202178 227338
rect 202346 227144 204110 227338
rect 204278 227144 205398 227338
rect 205566 227144 207330 227338
rect 207498 227144 209262 227338
rect 209430 227144 211194 227338
rect 211362 227144 212482 227338
rect 212650 227144 214414 227338
rect 214582 227144 216346 227338
rect 216514 227144 218278 227338
rect 218446 227144 219566 227338
rect 219734 227144 221498 227338
rect 221666 227144 223430 227338
rect 223598 227144 225362 227338
rect 225530 227144 226650 227338
rect 226818 227144 228582 227338
rect 228750 227144 230514 227338
rect 230682 227144 232446 227338
rect 232614 227144 233734 227338
rect 233902 227144 235666 227338
rect 235834 227144 237598 227338
rect 237766 227144 239530 227338
rect 239698 227144 240818 227338
rect 240986 227144 242750 227338
rect 242918 227144 244682 227338
rect 244850 227144 246614 227338
rect 246782 227144 247902 227338
rect 248070 227144 249834 227338
rect 250002 227144 251766 227338
rect 251934 227144 253698 227338
rect 253866 227144 254986 227338
rect 255154 227144 256918 227338
rect 257086 227144 258850 227338
rect 259018 227144 260782 227338
rect 260950 227144 262070 227338
rect 262238 227144 264002 227338
rect 264170 227144 265934 227338
rect 266102 227144 267866 227338
rect 268034 227144 269154 227338
rect 269322 227144 271086 227338
rect 271254 227144 273018 227338
rect 273186 227144 274950 227338
rect 275118 227144 276238 227338
rect 276406 227144 278170 227338
rect 278338 227144 280102 227338
rect 280270 227144 281390 227338
rect 281558 227144 283322 227338
rect 283490 227144 285254 227338
rect 285422 227144 287186 227338
rect 287354 227144 288474 227338
rect 288642 227144 290406 227338
rect 290574 227144 292338 227338
rect 292506 227144 294270 227338
rect 294438 227144 295558 227338
rect 295726 227144 297490 227338
rect 297658 227144 299422 227338
rect 299590 227144 301354 227338
rect 301522 227144 302642 227338
rect 302810 227144 304574 227338
rect 304742 227144 306506 227338
rect 306674 227144 308438 227338
rect 308606 227144 309726 227338
rect 309894 227144 311658 227338
rect 311826 227144 313590 227338
rect 313758 227144 315522 227338
rect 315690 227144 316810 227338
rect 316978 227144 318026 227338
rect 20 856 318026 227144
rect 130 734 1250 856
rect 1418 734 3182 856
rect 3350 734 5114 856
rect 5282 734 6402 856
rect 6570 734 8334 856
rect 8502 734 10266 856
rect 10434 734 12198 856
rect 12366 734 13486 856
rect 13654 734 15418 856
rect 15586 734 17350 856
rect 17518 734 19282 856
rect 19450 734 20570 856
rect 20738 734 22502 856
rect 22670 734 24434 856
rect 24602 734 26366 856
rect 26534 734 27654 856
rect 27822 734 29586 856
rect 29754 734 31518 856
rect 31686 734 33450 856
rect 33618 734 34738 856
rect 34906 734 36670 856
rect 36838 734 38602 856
rect 38770 734 40534 856
rect 40702 734 41822 856
rect 41990 734 43754 856
rect 43922 734 45686 856
rect 45854 734 47618 856
rect 47786 734 48906 856
rect 49074 734 50838 856
rect 51006 734 52770 856
rect 52938 734 54702 856
rect 54870 734 55990 856
rect 56158 734 57922 856
rect 58090 734 59854 856
rect 60022 734 61786 856
rect 61954 734 63074 856
rect 63242 734 65006 856
rect 65174 734 66938 856
rect 67106 734 68870 856
rect 69038 734 70158 856
rect 70326 734 72090 856
rect 72258 734 74022 856
rect 74190 734 75954 856
rect 76122 734 77242 856
rect 77410 734 79174 856
rect 79342 734 81106 856
rect 81274 734 82394 856
rect 82562 734 84326 856
rect 84494 734 86258 856
rect 86426 734 88190 856
rect 88358 734 89478 856
rect 89646 734 91410 856
rect 91578 734 93342 856
rect 93510 734 95274 856
rect 95442 734 96562 856
rect 96730 734 98494 856
rect 98662 734 100426 856
rect 100594 734 102358 856
rect 102526 734 103646 856
rect 103814 734 105578 856
rect 105746 734 107510 856
rect 107678 734 109442 856
rect 109610 734 110730 856
rect 110898 734 112662 856
rect 112830 734 114594 856
rect 114762 734 116526 856
rect 116694 734 117814 856
rect 117982 734 119746 856
rect 119914 734 121678 856
rect 121846 734 123610 856
rect 123778 734 124898 856
rect 125066 734 126830 856
rect 126998 734 128762 856
rect 128930 734 130694 856
rect 130862 734 131982 856
rect 132150 734 133914 856
rect 134082 734 135846 856
rect 136014 734 137778 856
rect 137946 734 139066 856
rect 139234 734 140998 856
rect 141166 734 142930 856
rect 143098 734 144862 856
rect 145030 734 146150 856
rect 146318 734 148082 856
rect 148250 734 150014 856
rect 150182 734 151946 856
rect 152114 734 153234 856
rect 153402 734 155166 856
rect 155334 734 157098 856
rect 157266 734 159030 856
rect 159198 734 160318 856
rect 160486 734 162250 856
rect 162418 734 164182 856
rect 164350 734 165470 856
rect 165638 734 167402 856
rect 167570 734 169334 856
rect 169502 734 171266 856
rect 171434 734 172554 856
rect 172722 734 174486 856
rect 174654 734 176418 856
rect 176586 734 178350 856
rect 178518 734 179638 856
rect 179806 734 181570 856
rect 181738 734 183502 856
rect 183670 734 185434 856
rect 185602 734 186722 856
rect 186890 734 188654 856
rect 188822 734 190586 856
rect 190754 734 192518 856
rect 192686 734 193806 856
rect 193974 734 195738 856
rect 195906 734 197670 856
rect 197838 734 199602 856
rect 199770 734 200890 856
rect 201058 734 202822 856
rect 202990 734 204754 856
rect 204922 734 206686 856
rect 206854 734 207974 856
rect 208142 734 209906 856
rect 210074 734 211838 856
rect 212006 734 213770 856
rect 213938 734 215058 856
rect 215226 734 216990 856
rect 217158 734 218922 856
rect 219090 734 220854 856
rect 221022 734 222142 856
rect 222310 734 224074 856
rect 224242 734 226006 856
rect 226174 734 227938 856
rect 228106 734 229226 856
rect 229394 734 231158 856
rect 231326 734 233090 856
rect 233258 734 235022 856
rect 235190 734 236310 856
rect 236478 734 238242 856
rect 238410 734 240174 856
rect 240342 734 242106 856
rect 242274 734 243394 856
rect 243562 734 245326 856
rect 245494 734 247258 856
rect 247426 734 248546 856
rect 248714 734 250478 856
rect 250646 734 252410 856
rect 252578 734 254342 856
rect 254510 734 255630 856
rect 255798 734 257562 856
rect 257730 734 259494 856
rect 259662 734 261426 856
rect 261594 734 262714 856
rect 262882 734 264646 856
rect 264814 734 266578 856
rect 266746 734 268510 856
rect 268678 734 269798 856
rect 269966 734 271730 856
rect 271898 734 273662 856
rect 273830 734 275594 856
rect 275762 734 276882 856
rect 277050 734 278814 856
rect 278982 734 280746 856
rect 280914 734 282678 856
rect 282846 734 283966 856
rect 284134 734 285898 856
rect 286066 734 287830 856
rect 287998 734 289762 856
rect 289930 734 291050 856
rect 291218 734 292982 856
rect 293150 734 294914 856
rect 295082 734 296846 856
rect 297014 734 298134 856
rect 298302 734 300066 856
rect 300234 734 301998 856
rect 302166 734 303930 856
rect 304098 734 305218 856
rect 305386 734 307150 856
rect 307318 734 309082 856
rect 309250 734 311014 856
rect 311182 734 312302 856
rect 312470 734 314234 856
rect 314402 734 316166 856
rect 316334 734 318026 856
<< metal3 >>
rect 0 227128 800 227248
rect 319200 227128 320000 227248
rect 0 225768 800 225888
rect 319200 225088 320000 225208
rect 0 223728 800 223848
rect 319200 223728 320000 223848
rect 0 221688 800 221808
rect 319200 221688 320000 221808
rect 0 219648 800 219768
rect 319200 219648 320000 219768
rect 0 218288 800 218408
rect 319200 217608 320000 217728
rect 0 216248 800 216368
rect 319200 216248 320000 216368
rect 0 214208 800 214328
rect 319200 214208 320000 214328
rect 0 212168 800 212288
rect 319200 212168 320000 212288
rect 0 210808 800 210928
rect 319200 210128 320000 210248
rect 0 208768 800 208888
rect 319200 208768 320000 208888
rect 0 206728 800 206848
rect 319200 206728 320000 206848
rect 0 204688 800 204808
rect 319200 204688 320000 204808
rect 0 203328 800 203448
rect 319200 202648 320000 202768
rect 0 201288 800 201408
rect 319200 201288 320000 201408
rect 0 199248 800 199368
rect 319200 199248 320000 199368
rect 0 197208 800 197328
rect 319200 197208 320000 197328
rect 0 195848 800 195968
rect 319200 195168 320000 195288
rect 0 193808 800 193928
rect 319200 193808 320000 193928
rect 0 191768 800 191888
rect 319200 191768 320000 191888
rect 0 189728 800 189848
rect 319200 189728 320000 189848
rect 0 188368 800 188488
rect 319200 187688 320000 187808
rect 0 186328 800 186448
rect 319200 186328 320000 186448
rect 0 184288 800 184408
rect 319200 184288 320000 184408
rect 0 182248 800 182368
rect 319200 182248 320000 182368
rect 0 180888 800 181008
rect 319200 180888 320000 181008
rect 0 178848 800 178968
rect 319200 178848 320000 178968
rect 0 176808 800 176928
rect 319200 176808 320000 176928
rect 0 174768 800 174888
rect 319200 174768 320000 174888
rect 0 173408 800 173528
rect 319200 173408 320000 173528
rect 0 171368 800 171488
rect 319200 171368 320000 171488
rect 0 169328 800 169448
rect 319200 169328 320000 169448
rect 0 167968 800 168088
rect 319200 167288 320000 167408
rect 0 165928 800 166048
rect 319200 165928 320000 166048
rect 0 163888 800 164008
rect 319200 163888 320000 164008
rect 0 161848 800 161968
rect 319200 161848 320000 161968
rect 0 160488 800 160608
rect 319200 159808 320000 159928
rect 0 158448 800 158568
rect 319200 158448 320000 158568
rect 0 156408 800 156528
rect 319200 156408 320000 156528
rect 0 154368 800 154488
rect 319200 154368 320000 154488
rect 0 153008 800 153128
rect 319200 152328 320000 152448
rect 0 150968 800 151088
rect 319200 150968 320000 151088
rect 0 148928 800 149048
rect 319200 148928 320000 149048
rect 0 146888 800 147008
rect 319200 146888 320000 147008
rect 0 145528 800 145648
rect 319200 144848 320000 144968
rect 0 143488 800 143608
rect 319200 143488 320000 143608
rect 0 141448 800 141568
rect 319200 141448 320000 141568
rect 0 139408 800 139528
rect 319200 139408 320000 139528
rect 0 138048 800 138168
rect 319200 137368 320000 137488
rect 0 136008 800 136128
rect 319200 136008 320000 136128
rect 0 133968 800 134088
rect 319200 133968 320000 134088
rect 0 131928 800 132048
rect 319200 131928 320000 132048
rect 0 130568 800 130688
rect 319200 129888 320000 130008
rect 0 128528 800 128648
rect 319200 128528 320000 128648
rect 0 126488 800 126608
rect 319200 126488 320000 126608
rect 0 124448 800 124568
rect 319200 124448 320000 124568
rect 0 123088 800 123208
rect 319200 122408 320000 122528
rect 0 121048 800 121168
rect 319200 121048 320000 121168
rect 0 119008 800 119128
rect 319200 119008 320000 119128
rect 0 116968 800 117088
rect 319200 116968 320000 117088
rect 0 115608 800 115728
rect 319200 114928 320000 115048
rect 0 113568 800 113688
rect 319200 113568 320000 113688
rect 0 111528 800 111648
rect 319200 111528 320000 111648
rect 0 109488 800 109608
rect 319200 109488 320000 109608
rect 0 108128 800 108248
rect 319200 107448 320000 107568
rect 0 106088 800 106208
rect 319200 106088 320000 106208
rect 0 104048 800 104168
rect 319200 104048 320000 104168
rect 0 102008 800 102128
rect 319200 102008 320000 102128
rect 0 100648 800 100768
rect 319200 99968 320000 100088
rect 0 98608 800 98728
rect 319200 98608 320000 98728
rect 0 96568 800 96688
rect 319200 96568 320000 96688
rect 0 94528 800 94648
rect 319200 94528 320000 94648
rect 0 93168 800 93288
rect 319200 93168 320000 93288
rect 0 91128 800 91248
rect 319200 91128 320000 91248
rect 0 89088 800 89208
rect 319200 89088 320000 89208
rect 0 87048 800 87168
rect 319200 87048 320000 87168
rect 0 85688 800 85808
rect 319200 85688 320000 85808
rect 0 83648 800 83768
rect 319200 83648 320000 83768
rect 0 81608 800 81728
rect 319200 81608 320000 81728
rect 0 80248 800 80368
rect 319200 79568 320000 79688
rect 0 78208 800 78328
rect 319200 78208 320000 78328
rect 0 76168 800 76288
rect 319200 76168 320000 76288
rect 0 74128 800 74248
rect 319200 74128 320000 74248
rect 0 72768 800 72888
rect 319200 72088 320000 72208
rect 0 70728 800 70848
rect 319200 70728 320000 70848
rect 0 68688 800 68808
rect 319200 68688 320000 68808
rect 0 66648 800 66768
rect 319200 66648 320000 66768
rect 0 65288 800 65408
rect 319200 64608 320000 64728
rect 0 63248 800 63368
rect 319200 63248 320000 63368
rect 0 61208 800 61328
rect 319200 61208 320000 61328
rect 0 59168 800 59288
rect 319200 59168 320000 59288
rect 0 57808 800 57928
rect 319200 57128 320000 57248
rect 0 55768 800 55888
rect 319200 55768 320000 55888
rect 0 53728 800 53848
rect 319200 53728 320000 53848
rect 0 51688 800 51808
rect 319200 51688 320000 51808
rect 0 50328 800 50448
rect 319200 49648 320000 49768
rect 0 48288 800 48408
rect 319200 48288 320000 48408
rect 0 46248 800 46368
rect 319200 46248 320000 46368
rect 0 44208 800 44328
rect 319200 44208 320000 44328
rect 0 42848 800 42968
rect 319200 42168 320000 42288
rect 0 40808 800 40928
rect 319200 40808 320000 40928
rect 0 38768 800 38888
rect 319200 38768 320000 38888
rect 0 36728 800 36848
rect 319200 36728 320000 36848
rect 0 35368 800 35488
rect 319200 34688 320000 34808
rect 0 33328 800 33448
rect 319200 33328 320000 33448
rect 0 31288 800 31408
rect 319200 31288 320000 31408
rect 0 29248 800 29368
rect 319200 29248 320000 29368
rect 0 27888 800 28008
rect 319200 27208 320000 27328
rect 0 25848 800 25968
rect 319200 25848 320000 25968
rect 0 23808 800 23928
rect 319200 23808 320000 23928
rect 0 21768 800 21888
rect 319200 21768 320000 21888
rect 0 20408 800 20528
rect 319200 19728 320000 19848
rect 0 18368 800 18488
rect 319200 18368 320000 18488
rect 0 16328 800 16448
rect 319200 16328 320000 16448
rect 0 14288 800 14408
rect 319200 14288 320000 14408
rect 0 12928 800 13048
rect 319200 12248 320000 12368
rect 0 10888 800 11008
rect 319200 10888 320000 11008
rect 0 8848 800 8968
rect 319200 8848 320000 8968
rect 0 6808 800 6928
rect 319200 6808 320000 6928
rect 0 5448 800 5568
rect 319200 5448 320000 5568
rect 0 3408 800 3528
rect 319200 3408 320000 3528
rect 0 1368 800 1488
rect 319200 1368 320000 1488
<< obsm3 >>
rect 880 227048 319120 227221
rect 800 225968 319200 227048
rect 880 225688 319200 225968
rect 800 225288 319200 225688
rect 800 225008 319120 225288
rect 800 223928 319200 225008
rect 880 223648 319120 223928
rect 800 221888 319200 223648
rect 880 221608 319120 221888
rect 800 219848 319200 221608
rect 880 219568 319120 219848
rect 800 218488 319200 219568
rect 880 218208 319200 218488
rect 800 217808 319200 218208
rect 800 217528 319120 217808
rect 800 216448 319200 217528
rect 880 216168 319120 216448
rect 800 214408 319200 216168
rect 880 214128 319120 214408
rect 800 212368 319200 214128
rect 880 212088 319120 212368
rect 800 211008 319200 212088
rect 880 210728 319200 211008
rect 800 210328 319200 210728
rect 800 210048 319120 210328
rect 800 208968 319200 210048
rect 880 208688 319120 208968
rect 800 206928 319200 208688
rect 880 206648 319120 206928
rect 800 204888 319200 206648
rect 880 204608 319120 204888
rect 800 203528 319200 204608
rect 880 203248 319200 203528
rect 800 202848 319200 203248
rect 800 202568 319120 202848
rect 800 201488 319200 202568
rect 880 201208 319120 201488
rect 800 199448 319200 201208
rect 880 199168 319120 199448
rect 800 197408 319200 199168
rect 880 197128 319120 197408
rect 800 196048 319200 197128
rect 880 195768 319200 196048
rect 800 195368 319200 195768
rect 800 195088 319120 195368
rect 800 194008 319200 195088
rect 880 193728 319120 194008
rect 800 191968 319200 193728
rect 880 191688 319120 191968
rect 800 189928 319200 191688
rect 880 189648 319120 189928
rect 800 188568 319200 189648
rect 880 188288 319200 188568
rect 800 187888 319200 188288
rect 800 187608 319120 187888
rect 800 186528 319200 187608
rect 880 186248 319120 186528
rect 800 184488 319200 186248
rect 880 184208 319120 184488
rect 800 182448 319200 184208
rect 880 182168 319120 182448
rect 800 181088 319200 182168
rect 880 180808 319120 181088
rect 800 179048 319200 180808
rect 880 178768 319120 179048
rect 800 177008 319200 178768
rect 880 176728 319120 177008
rect 800 174968 319200 176728
rect 880 174688 319120 174968
rect 800 173608 319200 174688
rect 880 173328 319120 173608
rect 800 171568 319200 173328
rect 880 171288 319120 171568
rect 800 169528 319200 171288
rect 880 169248 319120 169528
rect 800 168168 319200 169248
rect 880 167888 319200 168168
rect 800 167488 319200 167888
rect 800 167208 319120 167488
rect 800 166128 319200 167208
rect 880 165848 319120 166128
rect 800 164088 319200 165848
rect 880 163808 319120 164088
rect 800 162048 319200 163808
rect 880 161768 319120 162048
rect 800 160688 319200 161768
rect 880 160408 319200 160688
rect 800 160008 319200 160408
rect 800 159728 319120 160008
rect 800 158648 319200 159728
rect 880 158368 319120 158648
rect 800 156608 319200 158368
rect 880 156328 319120 156608
rect 800 154568 319200 156328
rect 880 154288 319120 154568
rect 800 153208 319200 154288
rect 880 152928 319200 153208
rect 800 152528 319200 152928
rect 800 152248 319120 152528
rect 800 151168 319200 152248
rect 880 150888 319120 151168
rect 800 149128 319200 150888
rect 880 148848 319120 149128
rect 800 147088 319200 148848
rect 880 146808 319120 147088
rect 800 145728 319200 146808
rect 880 145448 319200 145728
rect 800 145048 319200 145448
rect 800 144768 319120 145048
rect 800 143688 319200 144768
rect 880 143408 319120 143688
rect 800 141648 319200 143408
rect 880 141368 319120 141648
rect 800 139608 319200 141368
rect 880 139328 319120 139608
rect 800 138248 319200 139328
rect 880 137968 319200 138248
rect 800 137568 319200 137968
rect 800 137288 319120 137568
rect 800 136208 319200 137288
rect 880 135928 319120 136208
rect 800 134168 319200 135928
rect 880 133888 319120 134168
rect 800 132128 319200 133888
rect 880 131848 319120 132128
rect 800 130768 319200 131848
rect 880 130488 319200 130768
rect 800 130088 319200 130488
rect 800 129808 319120 130088
rect 800 128728 319200 129808
rect 880 128448 319120 128728
rect 800 126688 319200 128448
rect 880 126408 319120 126688
rect 800 124648 319200 126408
rect 880 124368 319120 124648
rect 800 123288 319200 124368
rect 880 123008 319200 123288
rect 800 122608 319200 123008
rect 800 122328 319120 122608
rect 800 121248 319200 122328
rect 880 120968 319120 121248
rect 800 119208 319200 120968
rect 880 118928 319120 119208
rect 800 117168 319200 118928
rect 880 116888 319120 117168
rect 800 115808 319200 116888
rect 880 115528 319200 115808
rect 800 115128 319200 115528
rect 800 114848 319120 115128
rect 800 113768 319200 114848
rect 880 113488 319120 113768
rect 800 111728 319200 113488
rect 880 111448 319120 111728
rect 800 109688 319200 111448
rect 880 109408 319120 109688
rect 800 108328 319200 109408
rect 880 108048 319200 108328
rect 800 107648 319200 108048
rect 800 107368 319120 107648
rect 800 106288 319200 107368
rect 880 106008 319120 106288
rect 800 104248 319200 106008
rect 880 103968 319120 104248
rect 800 102208 319200 103968
rect 880 101928 319120 102208
rect 800 100848 319200 101928
rect 880 100568 319200 100848
rect 800 100168 319200 100568
rect 800 99888 319120 100168
rect 800 98808 319200 99888
rect 880 98528 319120 98808
rect 800 96768 319200 98528
rect 880 96488 319120 96768
rect 800 94728 319200 96488
rect 880 94448 319120 94728
rect 800 93368 319200 94448
rect 880 93088 319120 93368
rect 800 91328 319200 93088
rect 880 91048 319120 91328
rect 800 89288 319200 91048
rect 880 89008 319120 89288
rect 800 87248 319200 89008
rect 880 86968 319120 87248
rect 800 85888 319200 86968
rect 880 85608 319120 85888
rect 800 83848 319200 85608
rect 880 83568 319120 83848
rect 800 81808 319200 83568
rect 880 81528 319120 81808
rect 800 80448 319200 81528
rect 880 80168 319200 80448
rect 800 79768 319200 80168
rect 800 79488 319120 79768
rect 800 78408 319200 79488
rect 880 78128 319120 78408
rect 800 76368 319200 78128
rect 880 76088 319120 76368
rect 800 74328 319200 76088
rect 880 74048 319120 74328
rect 800 72968 319200 74048
rect 880 72688 319200 72968
rect 800 72288 319200 72688
rect 800 72008 319120 72288
rect 800 70928 319200 72008
rect 880 70648 319120 70928
rect 800 68888 319200 70648
rect 880 68608 319120 68888
rect 800 66848 319200 68608
rect 880 66568 319120 66848
rect 800 65488 319200 66568
rect 880 65208 319200 65488
rect 800 64808 319200 65208
rect 800 64528 319120 64808
rect 800 63448 319200 64528
rect 880 63168 319120 63448
rect 800 61408 319200 63168
rect 880 61128 319120 61408
rect 800 59368 319200 61128
rect 880 59088 319120 59368
rect 800 58008 319200 59088
rect 880 57728 319200 58008
rect 800 57328 319200 57728
rect 800 57048 319120 57328
rect 800 55968 319200 57048
rect 880 55688 319120 55968
rect 800 53928 319200 55688
rect 880 53648 319120 53928
rect 800 51888 319200 53648
rect 880 51608 319120 51888
rect 800 50528 319200 51608
rect 880 50248 319200 50528
rect 800 49848 319200 50248
rect 800 49568 319120 49848
rect 800 48488 319200 49568
rect 880 48208 319120 48488
rect 800 46448 319200 48208
rect 880 46168 319120 46448
rect 800 44408 319200 46168
rect 880 44128 319120 44408
rect 800 43048 319200 44128
rect 880 42768 319200 43048
rect 800 42368 319200 42768
rect 800 42088 319120 42368
rect 800 41008 319200 42088
rect 880 40728 319120 41008
rect 800 38968 319200 40728
rect 880 38688 319120 38968
rect 800 36928 319200 38688
rect 880 36648 319120 36928
rect 800 35568 319200 36648
rect 880 35288 319200 35568
rect 800 34888 319200 35288
rect 800 34608 319120 34888
rect 800 33528 319200 34608
rect 880 33248 319120 33528
rect 800 31488 319200 33248
rect 880 31208 319120 31488
rect 800 29448 319200 31208
rect 880 29168 319120 29448
rect 800 28088 319200 29168
rect 880 27808 319200 28088
rect 800 27408 319200 27808
rect 800 27128 319120 27408
rect 800 26048 319200 27128
rect 880 25768 319120 26048
rect 800 24008 319200 25768
rect 880 23728 319120 24008
rect 800 21968 319200 23728
rect 880 21688 319120 21968
rect 800 20608 319200 21688
rect 880 20328 319200 20608
rect 800 19928 319200 20328
rect 800 19648 319120 19928
rect 800 18568 319200 19648
rect 880 18288 319120 18568
rect 800 16528 319200 18288
rect 880 16248 319120 16528
rect 800 14488 319200 16248
rect 880 14208 319120 14488
rect 800 13128 319200 14208
rect 880 12848 319200 13128
rect 800 12448 319200 12848
rect 800 12168 319120 12448
rect 800 11088 319200 12168
rect 880 10808 319120 11088
rect 800 9048 319200 10808
rect 880 8768 319120 9048
rect 800 7008 319200 8768
rect 880 6728 319120 7008
rect 800 5648 319200 6728
rect 880 5368 319120 5648
rect 800 3608 319200 5368
rect 880 3328 319120 3608
rect 800 2143 319200 3328
<< metal4 >>
rect 4208 2128 4528 225808
rect 14208 2128 14528 225808
rect 24208 2128 24528 225808
rect 34208 2128 34528 225808
rect 44208 205452 44528 225808
rect 54208 205452 54528 225808
rect 64208 205452 64528 225808
rect 74208 205452 74528 225808
rect 84208 205452 84528 225808
rect 94208 205452 94528 225808
rect 104208 205452 104528 225808
rect 114208 205452 114528 225808
rect 124208 205452 124528 225808
rect 134208 205452 134528 225808
rect 44208 101452 44528 122048
rect 54208 101452 54528 122048
rect 64208 101452 64528 122048
rect 74208 101452 74528 122048
rect 84208 101452 84528 122048
rect 94208 101452 94528 122048
rect 104208 101452 104528 122048
rect 114208 101452 114528 122048
rect 124208 101452 124528 122048
rect 134208 101452 134528 122048
rect 44208 2128 44528 18048
rect 54208 2128 54528 18048
rect 64208 2128 64528 18048
rect 74208 2128 74528 18048
rect 84208 2128 84528 18048
rect 94208 2128 94528 18048
rect 104208 2128 104528 18048
rect 114208 2128 114528 18048
rect 124208 2128 124528 18048
rect 134208 2128 134528 18048
rect 144208 2128 144528 225808
rect 154208 2128 154528 225808
rect 164208 2128 164528 225808
rect 174208 2128 174528 225808
rect 184208 205452 184528 225808
rect 194208 205452 194528 225808
rect 204208 205452 204528 225808
rect 214208 205452 214528 225808
rect 224208 205452 224528 225808
rect 234208 205452 234528 225808
rect 244208 205452 244528 225808
rect 254208 205452 254528 225808
rect 264208 205452 264528 225808
rect 274208 205452 274528 225808
rect 184208 101452 184528 122048
rect 194208 101452 194528 122048
rect 204208 101452 204528 122048
rect 214208 101452 214528 122048
rect 224208 101452 224528 122048
rect 234208 101452 234528 122048
rect 244208 101452 244528 122048
rect 254208 101452 254528 122048
rect 264208 101452 264528 122048
rect 274208 101452 274528 122048
rect 184208 2128 184528 18048
rect 194208 2128 194528 18048
rect 204208 2128 204528 18048
rect 214208 2128 214528 18048
rect 224208 2128 224528 18048
rect 234208 2128 234528 18048
rect 244208 2128 244528 18048
rect 254208 2128 254528 18048
rect 264208 2128 264528 18048
rect 274208 2128 274528 18048
rect 284208 2128 284528 225808
rect 294208 2128 294528 225808
rect 304208 2128 304528 225808
rect 314208 2128 314528 225808
<< obsm4 >>
rect 38883 205372 44128 207093
rect 44608 205372 54128 207093
rect 54608 205372 64128 207093
rect 64608 205372 74128 207093
rect 74608 205372 84128 207093
rect 84608 205372 94128 207093
rect 94608 205372 104128 207093
rect 104608 205372 114128 207093
rect 114608 205372 124128 207093
rect 124608 205372 134128 207093
rect 134608 205372 144128 207093
rect 38883 122128 144128 205372
rect 38883 101372 44128 122128
rect 44608 101372 54128 122128
rect 54608 101372 64128 122128
rect 64608 101372 74128 122128
rect 74608 101372 84128 122128
rect 84608 101372 94128 122128
rect 94608 101372 104128 122128
rect 104608 101372 114128 122128
rect 114608 101372 124128 122128
rect 124608 101372 134128 122128
rect 134608 101372 144128 122128
rect 38883 18128 144128 101372
rect 38883 16627 44128 18128
rect 44608 16627 54128 18128
rect 54608 16627 64128 18128
rect 64608 16627 74128 18128
rect 74608 16627 84128 18128
rect 84608 16627 94128 18128
rect 94608 16627 104128 18128
rect 104608 16627 114128 18128
rect 114608 16627 124128 18128
rect 124608 16627 134128 18128
rect 134608 16627 144128 18128
rect 144608 16627 154128 207093
rect 154608 16627 164128 207093
rect 164608 16627 174128 207093
rect 174608 205372 184128 207093
rect 184608 205372 194128 207093
rect 194608 205372 204128 207093
rect 204608 205372 214128 207093
rect 214608 205372 224128 207093
rect 224608 205372 234128 207093
rect 234608 205372 244128 207093
rect 244608 205372 254128 207093
rect 254608 205372 264128 207093
rect 264608 205372 274128 207093
rect 274608 205372 276677 207093
rect 174608 122128 276677 205372
rect 174608 101372 184128 122128
rect 184608 101372 194128 122128
rect 194608 101372 204128 122128
rect 204608 101372 214128 122128
rect 214608 101372 224128 122128
rect 224608 101372 234128 122128
rect 234608 101372 244128 122128
rect 244608 101372 254128 122128
rect 254608 101372 264128 122128
rect 264608 101372 274128 122128
rect 274608 101372 276677 122128
rect 174608 18128 276677 101372
rect 174608 16627 184128 18128
rect 184608 16627 194128 18128
rect 194608 16627 204128 18128
rect 204608 16627 214128 18128
rect 214608 16627 224128 18128
rect 224608 16627 234128 18128
rect 234608 16627 244128 18128
rect 244608 16627 254128 18128
rect 254608 16627 264128 18128
rect 264608 16627 274128 18128
rect 274608 16627 276677 18128
<< labels >>
rlabel metal2 s 262770 0 262826 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 319200 72088 320000 72208 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 138478 227200 138534 228000 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 319200 131928 320000 132048 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 124310 227200 124366 228000 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 319200 216248 320000 216368 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 147494 227200 147550 228000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 115294 227200 115350 228000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 129462 227200 129518 228000 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 319200 156408 320000 156528 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 57334 227200 57390 228000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 218334 227200 218390 228000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 121090 227200 121146 228000 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 170678 227200 170734 228000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 2594 227200 2650 228000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 232502 227200 232558 228000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 205454 227200 205510 228000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 319200 133968 320000 134088 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 304630 227200 304686 228000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 303986 0 304042 800 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 319200 113568 320000 113688 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 177762 227200 177818 228000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 182248 800 182368 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 319200 48288 320000 48408 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 319200 42168 320000 42288 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 209318 227200 209374 228000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 142342 227200 142398 228000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 94686 227200 94742 228000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 319200 49648 320000 49768 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 48318 227200 48374 228000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 53470 227200 53526 228000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 181626 0 181682 800 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 95974 227200 96030 228000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 233790 227200 233846 228000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 319200 63248 320000 63368 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 319200 225088 320000 225208 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 219648 800 219768 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 78586 227200 78642 228000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 212538 227200 212594 228000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 319200 154368 320000 154488 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 319200 189728 320000 189848 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 18694 227200 18750 228000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 81806 227200 81862 228000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 59266 227200 59322 228000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 97906 227200 97962 228000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 206728 800 206848 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 255042 227200 255098 228000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 242806 227200 242862 228000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 309782 227200 309838 228000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 0 199248 800 199368 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 74722 227200 74778 228000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 45098 227200 45154 228000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 302698 227200 302754 228000 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 319200 208768 320000 208888 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 319200 165928 320000 166048 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 319200 12248 320000 12368 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 319200 129888 320000 130008 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 319200 199248 320000 199368 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 319200 167288 320000 167408 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 41234 227200 41290 228000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 255686 0 255742 800 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 300122 0 300178 800 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 191768 800 191888 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 101770 227200 101826 228000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 269854 0 269910 800 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 319200 104048 320000 104168 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 308494 227200 308550 228000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 319200 195168 320000 195288 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 243450 0 243506 800 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 319200 159808 320000 159928 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 316866 227200 316922 228000 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 319200 137368 320000 137488 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 99838 227200 99894 228000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 296902 0 296958 800 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 319200 122408 320000 122528 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 184846 227200 184902 228000 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 157798 227200 157854 228000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 43166 227200 43222 228000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 319200 61208 320000 61328 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 262126 227200 262182 228000 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 319200 91128 320000 91248 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 319200 27208 320000 27328 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 166814 227200 166870 228000 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 90822 227200 90878 228000 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 319200 204688 320000 204808 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 319200 124448 320000 124568 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 195150 227200 195206 228000 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 319200 21768 320000 21888 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 240874 227200 240930 228000 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 218288 800 218408 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 319200 126488 320000 126608 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 221688 800 221808 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 312358 0 312414 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 247958 227200 248014 228000 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 156510 227200 156566 228000 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 265990 227200 266046 228000 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 319200 116968 320000 117088 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 203328 800 203448 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 230570 227200 230626 228000 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 261482 0 261538 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 60554 227200 60610 228000 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 273718 0 273774 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 71502 227200 71558 228000 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 319200 150968 320000 151088 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 319200 66648 320000 66768 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 319200 184288 320000 184408 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 253754 227200 253810 228000 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 52182 227200 52238 228000 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 319200 96568 320000 96688 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 319200 3408 320000 3528 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 186328 800 186448 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 319200 173408 320000 173528 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 319200 114928 320000 115048 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 213826 0 213882 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 145562 227200 145618 228000 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 171966 227200 172022 228000 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 5814 227200 5870 228000 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 260838 227200 260894 228000 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 311714 227200 311770 228000 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 319200 70728 320000 70848 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 319200 76168 320000 76288 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 319200 163888 320000 164008 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 136546 227200 136602 228000 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 239586 227200 239642 228000 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 50250 227200 50306 228000 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 306562 227200 306618 228000 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 319200 1368 320000 1488 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 273074 227200 273130 228000 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 67638 227200 67694 228000 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 319200 16328 320000 16448 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 319200 212168 320000 212288 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 34150 227200 34206 228000 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 159730 227200 159786 228000 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 319200 152328 320000 152448 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 319200 59168 320000 59288 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 319200 18368 320000 18488 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 319442 0 319498 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 114006 227200 114062 228000 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 319200 128528 320000 128648 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 319200 171368 320000 171488 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 319200 25848 320000 25968 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 319200 34688 320000 34808 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 319200 36728 320000 36848 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 275006 227200 275062 228000 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 154578 227200 154634 228000 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 319200 146888 320000 147008 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 140410 227200 140466 228000 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 110142 227200 110198 228000 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 204166 227200 204222 228000 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 55402 227200 55458 228000 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 16762 227200 16818 228000 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 319200 79568 320000 79688 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 299478 227200 299534 228000 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 14830 227200 14886 228000 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 319200 51688 320000 51808 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 319200 99968 320000 100088 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 108854 227200 108910 228000 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 223728 800 223848 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 188066 227200 188122 228000 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 211250 227200 211306 228000 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 246670 227200 246726 228000 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 294326 227200 294382 228000 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 161662 227200 161718 228000 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 319200 193808 320000 193928 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 319200 10888 320000 11008 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 278870 0 278926 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 92754 227200 92810 228000 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 297546 227200 297602 228000 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 225768 800 225888 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 169328 800 169448 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 319200 197208 320000 197328 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 319200 74128 320000 74248 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 319200 87048 320000 87168 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 264702 0 264758 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 69570 227200 69626 228000 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 316222 0 316278 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 66350 227200 66406 228000 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 319200 219648 320000 219768 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 225418 227200 225474 228000 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 319200 53728 320000 53848 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 198370 227200 198426 228000 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 319200 78208 320000 78328 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 30930 227200 30986 228000 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 309138 0 309194 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 104990 227200 105046 228000 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 202234 227200 202290 228000 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 287242 227200 287298 228000 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 210808 800 210928 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 264058 227200 264114 228000 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 319200 23808 320000 23928 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 150714 227200 150770 228000 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 131394 227200 131450 228000 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 122378 227200 122434 228000 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 276938 0 276994 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 315578 227200 315634 228000 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 143630 227200 143686 228000 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 214208 800 214328 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 319200 89088 320000 89208 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 319200 81608 320000 81728 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 301410 227200 301466 228000 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 256974 227200 257030 228000 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 179050 227200 179106 228000 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 211894 0 211950 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 11610 227200 11666 228000 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 319200 98608 320000 98728 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 319200 8848 320000 8968 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 292394 227200 292450 228000 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 152646 227200 152702 228000 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 36082 227200 36138 228000 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 182914 227200 182970 228000 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 294970 0 295026 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 254398 0 254454 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 319200 6808 320000 6928 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 28998 227200 29054 228000 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 106922 227200 106978 228000 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 87602 227200 87658 228000 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 268566 0 268622 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 319200 93168 320000 93288 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 197082 227200 197138 228000 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 189998 227200 190054 228000 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 191930 227200 191986 228000 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 202878 0 202934 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 278226 227200 278282 228000 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 135258 227200 135314 228000 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 163594 227200 163650 228000 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 209962 0 210018 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 73434 227200 73490 228000 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 271142 227200 271198 228000 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 319200 223728 320000 223848 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 7746 227200 7802 228000 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 276294 227200 276350 228000 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 319200 109488 320000 109608 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 173898 227200 173954 228000 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 313646 227200 313702 228000 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 319200 106088 320000 106208 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 226706 227200 226762 228000 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 258906 227200 258962 228000 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 319200 161848 320000 161968 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 207386 227200 207442 228000 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 319200 214208 320000 214328 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 319200 57128 320000 57248 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 319200 107448 320000 107568 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 319200 180888 320000 181008 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 319200 19728 320000 19848 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 319200 141448 320000 141568 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 318154 0 318210 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 311070 0 311126 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 319200 210128 320000 210248 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 319200 64608 320000 64728 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 285310 227200 285366 228000 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 319200 102008 320000 102128 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 318798 227200 318854 228000 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 288530 227200 288586 228000 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 126242 227200 126298 228000 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 80518 227200 80574 228000 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 319200 38768 320000 38888 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 319200 111528 320000 111648 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 319200 176808 320000 176928 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 295614 227200 295670 228000 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 12898 227200 12954 228000 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 62486 227200 62542 228000 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 9678 227200 9734 228000 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 319200 33328 320000 33448 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 319200 178848 320000 178968 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 175830 227200 175886 228000 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 133326 227200 133382 228000 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 319200 206728 320000 206848 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 208768 800 208888 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 117226 227200 117282 228000 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 319200 174768 320000 174888 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 237654 227200 237710 228000 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 32218 227200 32274 228000 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 267922 227200 267978 228000 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 281446 227200 281502 228000 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 283378 227200 283434 228000 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 193218 227200 193274 228000 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 319200 5448 320000 5568 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 39302 227200 39358 228000 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 186134 227200 186190 228000 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 662 227200 718 228000 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 319200 143488 320000 143608 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 319200 202648 320000 202768 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 201288 800 201408 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 302054 0 302110 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 319200 187688 320000 187808 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 149426 227200 149482 228000 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 319200 148928 320000 149048 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 319200 14288 320000 14408 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 128174 227200 128230 228000 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 25778 227200 25834 228000 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 319200 186328 320000 186448 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 284022 0 284078 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 46386 227200 46442 228000 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 216402 227200 216458 228000 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 38014 227200 38070 228000 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 64418 227200 64474 228000 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 44208 2128 44528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 64208 2128 64528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 84208 2128 84528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 104208 2128 104528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 124208 2128 124528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 184208 2128 184528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 204208 2128 204528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 224208 2128 224528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 244208 2128 244528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 264208 2128 264528 18048 6 vccd1
port 502 nsew power input
rlabel metal4 s 44208 101452 44528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 64208 101452 64528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 84208 101452 84528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 104208 101452 104528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 124208 101452 124528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 184208 101452 184528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 204208 101452 204528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 224208 101452 224528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 244208 101452 244528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 264208 101452 264528 122048 6 vccd1
port 502 nsew power input
rlabel metal4 s 4208 2128 4528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 24208 2128 24528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 44208 205452 44528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 64208 205452 64528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 84208 205452 84528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 104208 205452 104528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 124208 205452 124528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 144208 2128 144528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 164208 2128 164528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 184208 205452 184528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 204208 205452 204528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 224208 205452 224528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 244208 205452 244528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 264208 205452 264528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 284208 2128 284528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 304208 2128 304528 225808 6 vccd1
port 502 nsew power input
rlabel metal4 s 54208 2128 54528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 74208 2128 74528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 94208 2128 94528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 114208 2128 114528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 134208 2128 134528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 194208 2128 194528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 214208 2128 214528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234208 2128 234528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 254208 2128 254528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 274208 2128 274528 18048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 54208 101452 54528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 74208 101452 74528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 94208 101452 94528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 114208 101452 114528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 134208 101452 134528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 194208 101452 194528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 214208 101452 214528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234208 101452 234528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 254208 101452 254528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 274208 101452 274528 122048 6 vssd1
port 503 nsew ground input
rlabel metal4 s 14208 2128 14528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 34208 2128 34528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 54208 205452 54528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 74208 205452 74528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 94208 205452 94528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 114208 205452 114528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 134208 205452 134528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 154208 2128 154528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 174208 2128 174528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 194208 205452 194528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 214208 205452 214528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234208 205452 234528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 254208 205452 254528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 274208 205452 274528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 294208 2128 294528 225808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 314208 2128 314528 225808 6 vssd1
port 503 nsew ground input
rlabel metal3 s 319200 31288 320000 31408 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 21914 227200 21970 228000 6 wb_rst_i
port 505 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 164882 227200 164938 228000 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 103058 227200 103114 228000 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal3 s 0 216248 800 216368 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal3 s 319200 201288 320000 201408 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal3 s 319200 182248 320000 182368 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal3 s 319200 68688 320000 68808 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 168746 227200 168802 228000 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 251822 227200 251878 228000 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal3 s 319200 40808 320000 40928 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 19982 227200 20038 228000 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 85670 227200 85726 228000 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal3 s 319200 144848 320000 144968 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 290462 227200 290518 228000 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 219622 227200 219678 228000 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal3 s 319200 94528 320000 94648 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 214470 227200 214526 228000 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 285954 0 286010 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal3 s 319200 46248 320000 46368 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 88890 227200 88946 228000 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal3 s 319200 227128 320000 227248 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal3 s 319200 119008 320000 119128 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 200302 227200 200358 228000 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 269210 227200 269266 228000 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 23846 227200 23902 228000 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal3 s 319200 139408 320000 139528 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 280158 227200 280214 228000 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal3 s 319200 191768 320000 191888 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal3 s 319200 55768 320000 55888 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 249890 227200 249946 228000 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 83738 227200 83794 228000 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal3 s 319200 136008 320000 136128 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal3 s 319200 44208 320000 44328 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 289818 0 289874 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal3 s 319200 83648 320000 83768 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 244738 227200 244794 228000 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal3 s 319200 217608 320000 217728 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 291106 0 291162 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal3 s 319200 121048 320000 121168 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal3 s 319200 221688 320000 221808 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 235722 227200 235778 228000 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 217046 0 217102 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal3 s 0 227128 800 227248 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 112074 227200 112130 228000 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 180982 227200 181038 228000 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 119158 227200 119214 228000 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 228638 227200 228694 228000 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal3 s 319200 29248 320000 29368 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal3 s 0 174768 800 174888 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal3 s 319200 169328 320000 169448 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal3 s 319200 158448 320000 158568 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 223486 227200 223542 228000 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 221554 227200 221610 228000 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 27066 227200 27122 228000 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 76654 227200 76710 228000 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4526 227200 4582 228000 6 wbs_stb_i
port 608 nsew signal input
rlabel metal3 s 319200 85688 320000 85808 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 320000 228000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 25019978
string GDS_FILE /home/serdar/Desktop/openram_demo/openram_openmpw/openlane/openram_demo/runs/openram_demo/results/signoff/openram_demo.magic.gds
string GDS_START 10044160
<< end >>

