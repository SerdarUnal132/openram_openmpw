VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32_16_sky130
   CLASS BLOCK ;
   SIZE 347.18 BY 166.3 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.48 0.0 75.86 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.92 0.0 81.3 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.04 0.0 87.42 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  92.48 0.0 92.86 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.28 0.0 99.66 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.72 0.0 105.1 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.84 0.0 111.22 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.6 0.0 115.98 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.4 0.0 122.78 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.28 0.0 133.66 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.08 0.0 140.46 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.84 0.0 145.22 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 0.0 151.34 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  162.52 0.0 162.9 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.96 0.0 168.34 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.08 0.0 174.46 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  185.64 0.0 186.02 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 0.0 209.82 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.88 0.0 215.26 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 0.0 222.06 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 0.0 226.82 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.24 0.0 233.62 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 0.0 245.18 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 0.0 251.3 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 0.0 256.74 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  62.56 165.24 62.94 166.3 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  64.6 165.24 64.98 166.3 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  63.92 165.24 64.3 166.3 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  63.24 165.24 63.62 166.3 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  346.12 70.72 347.18 71.1 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  346.12 63.24 347.18 63.62 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.56 0.0 283.94 1.06 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 0.0 284.62 1.06 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 16.32 1.06 16.7 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  346.12 150.28 347.18 150.66 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 23.8 1.06 24.18 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  29.92 0.0 30.3 1.06 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 165.24 316.58 166.3 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  123.76 0.0 124.14 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  129.2 0.0 129.58 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  130.56 0.0 130.94 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  135.32 0.0 135.7 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.68 0.0 137.06 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.12 0.0 142.5 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.8 0.0 143.18 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 0.0 148.62 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.92 0.0 149.3 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  154.36 0.0 154.74 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.04 0.0 155.42 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 0.0 160.86 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 0.0 163.58 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 0.0 166.98 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.0 0.0 170.38 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  174.76 0.0 175.14 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.8 0.0 177.18 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 0.0 181.26 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 0.0 186.7 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  188.36 0.0 188.74 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 0.0 192.14 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 0.0 198.26 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.24 0.0 199.62 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 0.0 210.5 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 0.0 211.86 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 0.0 217.3 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 0.0 223.42 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  123.76 165.24 124.14 166.3 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  129.2 165.24 129.58 166.3 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  130.56 165.24 130.94 166.3 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  135.32 165.24 135.7 166.3 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.68 165.24 137.06 166.3 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.12 165.24 142.5 166.3 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 165.24 143.86 166.3 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.56 165.24 147.94 166.3 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  149.6 165.24 149.98 166.3 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  154.36 165.24 154.74 166.3 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.72 165.24 156.1 166.3 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 165.24 160.86 166.3 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 165.24 162.22 166.3 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 165.24 166.98 166.3 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.96 165.24 168.34 166.3 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 165.24 173.78 166.3 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  174.08 165.24 174.46 166.3 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 165.24 179.22 166.3 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 165.24 180.58 166.3 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 165.24 185.34 166.3 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 165.24 186.7 166.3 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 165.24 192.14 166.3 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 165.24 193.5 166.3 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 165.24 198.26 166.3 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.24 165.24 199.62 166.3 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 165.24 204.38 166.3 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 165.24 205.74 166.3 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.8 165.24 211.18 166.3 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 165.24 211.86 166.3 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 165.24 217.3 166.3 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 165.24 217.98 166.3 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 165.24 223.42 166.3 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  340.68 4.76 342.42 161.54 ;
         LAYER met3 ;
         RECT  4.76 4.76 342.42 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 161.54 ;
         LAYER met3 ;
         RECT  4.76 159.8 342.42 161.54 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  1.36 1.36 345.82 3.1 ;
         LAYER met3 ;
         RECT  1.36 163.2 345.82 164.94 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 164.94 ;
         LAYER met4 ;
         RECT  344.08 1.36 345.82 164.94 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 346.56 165.68 ;
   LAYER  met2 ;
      RECT  0.62 0.62 346.56 165.68 ;
   LAYER  met3 ;
      RECT  0.62 70.12 345.52 71.7 ;
      RECT  345.52 64.22 346.56 70.12 ;
      RECT  1.66 15.72 345.52 17.3 ;
      RECT  1.66 17.3 345.52 70.12 ;
      RECT  345.52 71.7 346.56 149.68 ;
      RECT  0.62 17.3 1.66 23.2 ;
      RECT  0.62 24.78 1.66 70.12 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 15.72 ;
      RECT  4.16 7.1 343.02 15.72 ;
      RECT  343.02 4.16 345.52 7.1 ;
      RECT  343.02 7.1 345.52 15.72 ;
      RECT  0.62 71.7 4.16 159.2 ;
      RECT  0.62 159.2 4.16 162.14 ;
      RECT  4.16 71.7 343.02 159.2 ;
      RECT  343.02 71.7 345.52 159.2 ;
      RECT  343.02 159.2 345.52 162.14 ;
      RECT  345.52 0.62 346.42 0.76 ;
      RECT  345.52 3.7 346.42 62.64 ;
      RECT  346.42 0.62 346.56 0.76 ;
      RECT  346.42 0.76 346.56 3.7 ;
      RECT  346.42 3.7 346.56 62.64 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 15.72 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 15.72 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 343.02 0.76 ;
      RECT  4.16 3.7 343.02 4.16 ;
      RECT  343.02 0.62 345.52 0.76 ;
      RECT  343.02 3.7 345.52 4.16 ;
      RECT  345.52 151.26 346.42 162.6 ;
      RECT  345.52 165.54 346.42 165.68 ;
      RECT  346.42 151.26 346.56 162.6 ;
      RECT  346.42 162.6 346.56 165.54 ;
      RECT  346.42 165.54 346.56 165.68 ;
      RECT  0.62 162.14 0.76 162.6 ;
      RECT  0.62 162.6 0.76 165.54 ;
      RECT  0.62 165.54 0.76 165.68 ;
      RECT  0.76 162.14 4.16 162.6 ;
      RECT  0.76 165.54 4.16 165.68 ;
      RECT  4.16 162.14 343.02 162.6 ;
      RECT  4.16 165.54 343.02 165.68 ;
      RECT  343.02 162.14 345.52 162.6 ;
      RECT  343.02 165.54 345.52 165.68 ;
   LAYER  met4 ;
      RECT  74.88 1.66 76.46 165.68 ;
      RECT  76.46 0.62 80.32 1.66 ;
      RECT  81.9 0.62 86.44 1.66 ;
      RECT  88.02 0.62 91.88 1.66 ;
      RECT  93.46 0.62 98.68 1.66 ;
      RECT  100.26 0.62 104.12 1.66 ;
      RECT  105.7 0.62 110.24 1.66 ;
      RECT  111.82 0.62 115.0 1.66 ;
      RECT  116.58 0.62 121.8 1.66 ;
      RECT  227.42 0.62 232.64 1.66 ;
      RECT  234.22 0.62 238.76 1.66 ;
      RECT  240.34 0.62 244.2 1.66 ;
      RECT  245.78 0.62 250.32 1.66 ;
      RECT  251.9 0.62 255.76 1.66 ;
      RECT  61.96 1.66 63.54 164.64 ;
      RECT  63.54 1.66 74.88 164.64 ;
      RECT  65.58 164.64 74.88 165.68 ;
      RECT  257.34 0.62 282.96 1.66 ;
      RECT  30.9 0.62 74.88 1.66 ;
      RECT  76.46 1.66 315.6 164.64 ;
      RECT  315.6 1.66 317.18 164.64 ;
      RECT  124.74 0.62 126.56 1.66 ;
      RECT  128.14 0.62 128.6 1.66 ;
      RECT  131.54 0.62 132.68 1.66 ;
      RECT  134.26 0.62 134.72 1.66 ;
      RECT  137.66 0.62 139.48 1.66 ;
      RECT  141.06 0.62 141.52 1.66 ;
      RECT  143.78 0.62 144.24 1.66 ;
      RECT  145.82 0.62 147.64 1.66 ;
      RECT  149.9 0.62 150.36 1.66 ;
      RECT  151.94 0.62 153.76 1.66 ;
      RECT  157.38 0.62 159.88 1.66 ;
      RECT  161.46 0.62 161.92 1.66 ;
      RECT  164.18 0.62 166.0 1.66 ;
      RECT  168.94 0.62 169.4 1.66 ;
      RECT  170.98 0.62 172.12 1.66 ;
      RECT  175.74 0.62 176.2 1.66 ;
      RECT  177.78 0.62 179.6 1.66 ;
      RECT  181.86 0.62 185.04 1.66 ;
      RECT  187.3 0.62 187.76 1.66 ;
      RECT  189.34 0.62 191.16 1.66 ;
      RECT  194.1 0.62 196.6 1.66 ;
      RECT  200.22 0.62 202.72 1.66 ;
      RECT  206.34 0.62 208.84 1.66 ;
      RECT  212.46 0.62 214.28 1.66 ;
      RECT  215.86 0.62 216.32 1.66 ;
      RECT  218.58 0.62 221.08 1.66 ;
      RECT  224.02 0.62 225.84 1.66 ;
      RECT  76.46 164.64 123.16 165.68 ;
      RECT  124.74 164.64 128.6 165.68 ;
      RECT  131.54 164.64 134.72 165.68 ;
      RECT  137.66 164.64 141.52 165.68 ;
      RECT  144.46 164.64 146.96 165.68 ;
      RECT  148.54 164.64 149.0 165.68 ;
      RECT  150.58 164.64 153.76 165.68 ;
      RECT  156.7 164.64 159.88 165.68 ;
      RECT  162.82 164.64 166.0 165.68 ;
      RECT  168.94 164.64 172.8 165.68 ;
      RECT  175.06 164.64 178.24 165.68 ;
      RECT  181.18 164.64 184.36 165.68 ;
      RECT  187.3 164.64 191.16 165.68 ;
      RECT  194.1 164.64 197.28 165.68 ;
      RECT  200.22 164.64 203.4 165.68 ;
      RECT  206.34 164.64 210.2 165.68 ;
      RECT  212.46 164.64 216.32 165.68 ;
      RECT  218.58 164.64 222.44 165.68 ;
      RECT  224.02 164.64 315.6 165.68 ;
      RECT  317.18 1.66 340.08 4.16 ;
      RECT  317.18 4.16 340.08 162.14 ;
      RECT  317.18 162.14 340.08 164.64 ;
      RECT  340.08 1.66 343.02 4.16 ;
      RECT  340.08 162.14 343.02 164.64 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 162.14 7.1 164.64 ;
      RECT  7.1 1.66 61.96 4.16 ;
      RECT  7.1 4.16 61.96 162.14 ;
      RECT  7.1 162.14 61.96 164.64 ;
      RECT  0.62 164.64 0.76 165.54 ;
      RECT  0.62 165.54 0.76 165.68 ;
      RECT  0.76 165.54 3.7 165.68 ;
      RECT  3.7 164.64 61.96 165.54 ;
      RECT  3.7 165.54 61.96 165.68 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 29.32 0.76 ;
      RECT  3.7 0.76 29.32 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 162.14 ;
      RECT  3.7 4.16 4.16 162.14 ;
      RECT  0.62 162.14 0.76 164.64 ;
      RECT  3.7 162.14 4.16 164.64 ;
      RECT  285.22 0.62 343.48 0.76 ;
      RECT  285.22 0.76 343.48 1.66 ;
      RECT  343.48 0.62 346.42 0.76 ;
      RECT  346.42 0.62 346.56 0.76 ;
      RECT  346.42 0.76 346.56 1.66 ;
      RECT  317.18 164.64 343.48 165.54 ;
      RECT  317.18 165.54 343.48 165.68 ;
      RECT  343.48 165.54 346.42 165.68 ;
      RECT  346.42 164.64 346.56 165.54 ;
      RECT  346.42 165.54 346.56 165.68 ;
      RECT  343.02 1.66 343.48 4.16 ;
      RECT  346.42 1.66 346.56 4.16 ;
      RECT  343.02 4.16 343.48 162.14 ;
      RECT  346.42 4.16 346.56 162.14 ;
      RECT  343.02 162.14 343.48 164.64 ;
      RECT  346.42 162.14 346.56 164.64 ;
   END
END    sram_32_16_sky130
END    LIBRARY
